`define toAscii(x) { x / 8'ha + 8'h30, x % 8'ha + 8'h30 }

module RocketTile(
`ifdef MULTICORE
  input         cov_store,
  input         cov_restore,
  input [7:0]   proc_num,
`endif
  input         clock,
  input         reset,
  input         auto_intsink_in_sync_0,
  input         auto_int_in_xing_in_2_sync_0,
  input         auto_int_in_xing_in_1_sync_0,
  input         auto_int_in_xing_in_0_sync_0,
  input         auto_int_in_xing_in_0_sync_1,
  input         auto_tl_master_xing_out_a_ready,
  output        auto_tl_master_xing_out_a_valid,
  output [2:0]  auto_tl_master_xing_out_a_bits_opcode,
  output [2:0]  auto_tl_master_xing_out_a_bits_param,
  output [3:0]  auto_tl_master_xing_out_a_bits_size,
  output [1:0]  auto_tl_master_xing_out_a_bits_source,
  output [31:0] auto_tl_master_xing_out_a_bits_address,
  output [7:0]  auto_tl_master_xing_out_a_bits_mask,
  output [63:0] auto_tl_master_xing_out_a_bits_data,
  output        auto_tl_master_xing_out_a_bits_corrupt,
  output        auto_tl_master_xing_out_b_ready,
  input         auto_tl_master_xing_out_b_valid,
  input  [2:0]  auto_tl_master_xing_out_b_bits_opcode,
  input  [1:0]  auto_tl_master_xing_out_b_bits_param,
  input  [3:0]  auto_tl_master_xing_out_b_bits_size,
  input  [1:0]  auto_tl_master_xing_out_b_bits_source,
  input  [31:0] auto_tl_master_xing_out_b_bits_address,
  input  [7:0]  auto_tl_master_xing_out_b_bits_mask,
  input  [63:0] auto_tl_master_xing_out_b_bits_data,
  input         auto_tl_master_xing_out_b_bits_corrupt,
  input         auto_tl_master_xing_out_c_ready,
  output        auto_tl_master_xing_out_c_valid,
  output [2:0]  auto_tl_master_xing_out_c_bits_opcode,
  output [2:0]  auto_tl_master_xing_out_c_bits_param,
  output [3:0]  auto_tl_master_xing_out_c_bits_size,
  output [1:0]  auto_tl_master_xing_out_c_bits_source,
  output [31:0] auto_tl_master_xing_out_c_bits_address,
  output [63:0] auto_tl_master_xing_out_c_bits_data,
  output        auto_tl_master_xing_out_c_bits_corrupt,
  output        auto_tl_master_xing_out_d_ready,
  input         auto_tl_master_xing_out_d_valid,
  input  [2:0]  auto_tl_master_xing_out_d_bits_opcode,
  input  [1:0]  auto_tl_master_xing_out_d_bits_param,
  input  [3:0]  auto_tl_master_xing_out_d_bits_size,
  input  [1:0]  auto_tl_master_xing_out_d_bits_source,
  input  [1:0]  auto_tl_master_xing_out_d_bits_sink,
  input         auto_tl_master_xing_out_d_bits_denied,
  input  [63:0] auto_tl_master_xing_out_d_bits_data,
  input         auto_tl_master_xing_out_d_bits_corrupt,
  input         auto_tl_master_xing_out_e_ready,
  output        auto_tl_master_xing_out_e_valid,
  output [1:0]  auto_tl_master_xing_out_e_bits_sink,
  output        auto_wfi_out_0,
  output        auto_cease_out_0,
  output        auto_halt_out_0,
  input  [31:0] auto_reset_vector_in,
  input         auto_hartid_in,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         ptw_halt,
  input         resetVectorNode_halt,
  input         dcacheArb_halt,
  input         tlMasterXbar_halt,
  input         dcache_halt,
  input         intsink_3_halt,
  input         intsink_1_halt,
  input         buffer_halt,
  input         core_halt,
  input         fpuOpt_halt,
  input         intXbar_halt,
  input         frontend_halt,
  input         hartIdNode_halt,
  input         intsink_halt,
  input         intsink_2_halt,
  output [19:0] FPU_regstate,		//Jaewon_FPU_regstate
    output [29:0] FPU_covSum,		//Jaewon_FPU_covSum
    output [19:0] PTW_regstate,			//Jaewon_PTW_regstate
    output [29:0] PTW_covSum,			//Jaewon_PTW_covSum
    output [19:0] DCache_regstate,		//Jaewon_DCache_regstate
    output [29:0] DCache_covSum,		//Jaewon_DCache_covSum
    output [5:0]	 Frontend_regstate,	//Jaewon_Frontend_regstate
    output [29:0] Frontend_covSum,		//Jaewon_Frontend_covSum
    output [63:0] Frontend_covmap,		//Jaewon_Frontend_covmap
    output [19:0] Rocket_regstate,			//Jaewon_Rocket_regstate
    output [29:0] Rocket_covSum				//Jaewon_Rocket_covSum
);

  reg debug_print;
  initial begin
    if (!$value$plusargs("DEBUG=%d", debug_print)) begin
      debug_print = 0;
    end
  end

  always @(posedge clock) begin
    if (debug_print) begin
      if (core.coreMonitorBundle_valid & ~core.reset) begin
        $fwrite(32'h80000001, "%d 0x%x ", core.io_hartid, core.coreMonitorBundle_pc);
        $fwrite(32'h80000001,"(0x%x) DASM(%x)\n", core.coreMonitorBundle_inst, core.coreMonitorBundle_inst); // @[core.scala 1258:17]
      end
    end
  end

`ifdef MULTICORE
  integer i;
  integer fd;
  integer c;
  reg [8*100:1] out;
  initial begin
    if ($value$plusargs("OUT=%s", out)) begin
      $display("Output directory: %0s\n", out);
    end
  end
  always @(posedge clock) begin
    if (cov_restore) begin
      fd = $fopen({out, "/covmap/ptw.PTW_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "ptw.PTW_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          ptw.PTW_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/dcacheArb.HellaCacheArbiter_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "dcacheArb.HellaCacheArbiter_cov");
      else begin
        for (i=0; i<2; i=i+1) begin
          c = $fgetc(fd);
          dcacheArb.HellaCacheArbiter_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/tlMasterXbar.TLXbar_7_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "tlMasterXbar.TLXbar_7_cov");
      else begin
        for (i=0; i<8; i=i+1) begin
          c = $fgetc(fd);
          tlMasterXbar.TLXbar_7_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/dcache.DCache_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "dcache.DCache_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          dcache.DCache_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/dcache.pma_checker.TLB_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "dcache.pma_checker.TLB_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          dcache.pma_checker.TLB_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/dcache.tlb.TLB_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "dcache.tlb.TLB_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          dcache.tlb.TLB_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/core.Rocket_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "core.Rocket_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          core.Rocket_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/core.csr.CSRFile_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "core.csr.CSRFile_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          core.csr.CSRFile_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/core.div.MulDiv_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "core.div.MulDiv_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          core.div.MulDiv_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/core.ibuf.IBuf_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "core.ibuf.IBuf_cov");
      else begin
        for (i=0; i<4; i=i+1) begin
          c = $fgetc(fd);
          core.ibuf.IBuf_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.FPU_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.FPU_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.FPU_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.divSqrt_1.divSqrtRecFNToRaw.divSqrtRawFN.DivSqrtRawFN_small_1_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.divSqrt_1.divSqrtRecFNToRaw.divSqrtRawFN.DivSqrtRawFN_small_1_cov");
      else begin
        for (i=0; i<32; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.divSqrt_1.divSqrtRecFNToRaw.divSqrtRawFN.DivSqrtRawFN_small_1_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.ifpu.IntToFP_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.ifpu.IntToFP_cov");
      else begin
        for (i=0; i<32; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.ifpu.IntToFP_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.divSqrt.divSqrtRecFNToRaw.divSqrtRawFN.DivSqrtRawFN_small_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.divSqrt.divSqrtRecFNToRaw.divSqrtRawFN.DivSqrtRawFN_small_cov");
      else begin
        for (i=0; i<32; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.divSqrt.divSqrtRecFNToRaw.divSqrtRawFN.DivSqrtRawFN_small_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.fpmu.FPToFP_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.fpmu.FPToFP_cov");
      else begin
        for (i=0; i<128; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.fpmu.FPToFP_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.dfma.fma.MulAddRecFNPipe_1_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.dfma.fma.MulAddRecFNPipe_1_cov");
      else begin
        for (i=0; i<2; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.dfma.fma.MulAddRecFNPipe_1_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.fpiu.FPToInt_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.fpiu.FPToInt_cov");
      else begin
        for (i=0; i<32; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.fpiu.FPToInt_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.sfma.fma.MulAddRecFNPipe_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.sfma.fma.MulAddRecFNPipe_cov");
      else begin
        for (i=0; i<2; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.sfma.fma.MulAddRecFNPipe_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/frontend.Frontend_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "frontend.Frontend_cov");
      else begin
        for (i=0; i<64; i=i+1) begin
          c = $fgetc(fd);
          frontend.Frontend_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/frontend.icache.ICache_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "frontend.icache.ICache_cov");
      else begin
        for (i=0; i<64; i=i+1) begin
          c = $fgetc(fd);
          frontend.icache.ICache_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/frontend.fq.ShiftQueue_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "frontend.fq.ShiftQueue_cov");
      else begin
        for (i=0; i<2; i=i+1) begin
          c = $fgetc(fd);
          frontend.fq.ShiftQueue_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/frontend.tlb.TLB_1_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "frontend.tlb.TLB_1_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          frontend.tlb.TLB_1_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/frontend.btb.BTB_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "frontend.btb.BTB_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          frontend.btb.BTB_cov[i] = c[0];
        end
        $fclose(fd);
      end
    end
    if (cov_store) begin
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/ptw.PTW_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", ptw.PTW_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/dcacheArb.HellaCacheArbiter_cov.dat"}, "w");
      for (i=0; i<2; i=i+1)
        $fwrite(fd, "%0b", dcacheArb.HellaCacheArbiter_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/tlMasterXbar.TLXbar_7_cov.dat"}, "w");
      for (i=0; i<8; i=i+1)
        $fwrite(fd, "%0b", tlMasterXbar.TLXbar_7_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/dcache.DCache_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", dcache.DCache_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/dcache.pma_checker.TLB_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", dcache.pma_checker.TLB_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/dcache.tlb.TLB_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", dcache.tlb.TLB_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/core.Rocket_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", core.Rocket_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/core.csr.CSRFile_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", core.csr.CSRFile_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/core.div.MulDiv_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", core.div.MulDiv_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/core.ibuf.IBuf_cov.dat"}, "w");
      for (i=0; i<4; i=i+1)
        $fwrite(fd, "%0b", core.ibuf.IBuf_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/fpuOpt.FPU_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.FPU_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/fpuOpt.divSqrt_1.divSqrtRecFNToRaw.divSqrtRawFN.DivSqrtRawFN_small_1_cov.dat"}, "w");
      for (i=0; i<32; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.divSqrt_1.divSqrtRecFNToRaw.divSqrtRawFN.DivSqrtRawFN_small_1_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/fpuOpt.ifpu.IntToFP_cov.dat"}, "w");
      for (i=0; i<32; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.ifpu.IntToFP_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/fpuOpt.divSqrt.divSqrtRecFNToRaw.divSqrtRawFN.DivSqrtRawFN_small_cov.dat"}, "w");
      for (i=0; i<32; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.divSqrt.divSqrtRecFNToRaw.divSqrtRawFN.DivSqrtRawFN_small_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/fpuOpt.fpmu.FPToFP_cov.dat"}, "w");
      for (i=0; i<128; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.fpmu.FPToFP_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/fpuOpt.dfma.fma.MulAddRecFNPipe_1_cov.dat"}, "w");
      for (i=0; i<2; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.dfma.fma.MulAddRecFNPipe_1_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/fpuOpt.fpiu.FPToInt_cov.dat"}, "w");
      for (i=0; i<32; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.fpiu.FPToInt_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/fpuOpt.sfma.fma.MulAddRecFNPipe_cov.dat"}, "w");
      for (i=0; i<2; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.sfma.fma.MulAddRecFNPipe_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/frontend.Frontend_cov.dat"}, "w");
      for (i=0; i<64; i=i+1)
        $fwrite(fd, "%0b", frontend.Frontend_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/frontend.icache.ICache_cov.dat"}, "w");
      for (i=0; i<64; i=i+1)
        $fwrite(fd, "%0b", frontend.icache.ICache_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/frontend.fq.ShiftQueue_cov.dat"}, "w");
      for (i=0; i<2; i=i+1)
        $fwrite(fd, "%0b", frontend.fq.ShiftQueue_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/frontend.tlb.TLB_1_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", frontend.tlb.TLB_1_cov[i]);
      $fclose(fd);
      fd = $fopen({{{out, "/covmap-"}, `toAscii(proc_num)}, "/frontend.btb.BTB_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", frontend.btb.BTB_cov[i]);
      $fclose(fd);
    end
  end
`endif
  wire  tlMasterXbar_clock; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_reset; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_1_a_ready; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_1_a_valid; // @[BaseTile.scala 190:42]
  wire [31:0] tlMasterXbar_auto_in_1_a_bits_address; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_1_d_valid; // @[BaseTile.scala 190:42]
  wire [2:0] tlMasterXbar_auto_in_1_d_bits_opcode; // @[BaseTile.scala 190:42]
  wire [3:0] tlMasterXbar_auto_in_1_d_bits_size; // @[BaseTile.scala 190:42]
  wire [63:0] tlMasterXbar_auto_in_1_d_bits_data; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_1_d_bits_corrupt; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_a_ready; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_a_valid; // @[BaseTile.scala 190:42]
  wire [2:0] tlMasterXbar_auto_in_0_a_bits_opcode; // @[BaseTile.scala 190:42]
  wire [2:0] tlMasterXbar_auto_in_0_a_bits_param; // @[BaseTile.scala 190:42]
  wire [3:0] tlMasterXbar_auto_in_0_a_bits_size; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_a_bits_source; // @[BaseTile.scala 190:42]
  wire [31:0] tlMasterXbar_auto_in_0_a_bits_address; // @[BaseTile.scala 190:42]
  wire [7:0] tlMasterXbar_auto_in_0_a_bits_mask; // @[BaseTile.scala 190:42]
  wire [63:0] tlMasterXbar_auto_in_0_a_bits_data; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_b_ready; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_b_valid; // @[BaseTile.scala 190:42]
  wire [1:0] tlMasterXbar_auto_in_0_b_bits_param; // @[BaseTile.scala 190:42]
  wire [3:0] tlMasterXbar_auto_in_0_b_bits_size; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_b_bits_source; // @[BaseTile.scala 190:42]
  wire [31:0] tlMasterXbar_auto_in_0_b_bits_address; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_c_ready; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_c_valid; // @[BaseTile.scala 190:42]
  wire [2:0] tlMasterXbar_auto_in_0_c_bits_opcode; // @[BaseTile.scala 190:42]
  wire [2:0] tlMasterXbar_auto_in_0_c_bits_param; // @[BaseTile.scala 190:42]
  wire [3:0] tlMasterXbar_auto_in_0_c_bits_size; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_c_bits_source; // @[BaseTile.scala 190:42]
  wire [31:0] tlMasterXbar_auto_in_0_c_bits_address; // @[BaseTile.scala 190:42]
  wire [63:0] tlMasterXbar_auto_in_0_c_bits_data; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_d_ready; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_d_valid; // @[BaseTile.scala 190:42]
  wire [2:0] tlMasterXbar_auto_in_0_d_bits_opcode; // @[BaseTile.scala 190:42]
  wire [1:0] tlMasterXbar_auto_in_0_d_bits_param; // @[BaseTile.scala 190:42]
  wire [3:0] tlMasterXbar_auto_in_0_d_bits_size; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_d_bits_source; // @[BaseTile.scala 190:42]
  wire [1:0] tlMasterXbar_auto_in_0_d_bits_sink; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_d_bits_denied; // @[BaseTile.scala 190:42]
  wire [63:0] tlMasterXbar_auto_in_0_d_bits_data; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_e_ready; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_in_0_e_valid; // @[BaseTile.scala 190:42]
  wire [1:0] tlMasterXbar_auto_in_0_e_bits_sink; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_a_ready; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_a_valid; // @[BaseTile.scala 190:42]
  wire [2:0] tlMasterXbar_auto_out_a_bits_opcode; // @[BaseTile.scala 190:42]
  wire [2:0] tlMasterXbar_auto_out_a_bits_param; // @[BaseTile.scala 190:42]
  wire [3:0] tlMasterXbar_auto_out_a_bits_size; // @[BaseTile.scala 190:42]
  wire [1:0] tlMasterXbar_auto_out_a_bits_source; // @[BaseTile.scala 190:42]
  wire [31:0] tlMasterXbar_auto_out_a_bits_address; // @[BaseTile.scala 190:42]
  wire [7:0] tlMasterXbar_auto_out_a_bits_mask; // @[BaseTile.scala 190:42]
  wire [63:0] tlMasterXbar_auto_out_a_bits_data; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_a_bits_corrupt; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_b_ready; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_b_valid; // @[BaseTile.scala 190:42]
  wire [2:0] tlMasterXbar_auto_out_b_bits_opcode; // @[BaseTile.scala 190:42]
  wire [1:0] tlMasterXbar_auto_out_b_bits_param; // @[BaseTile.scala 190:42]
  wire [3:0] tlMasterXbar_auto_out_b_bits_size; // @[BaseTile.scala 190:42]
  wire [1:0] tlMasterXbar_auto_out_b_bits_source; // @[BaseTile.scala 190:42]
  wire [31:0] tlMasterXbar_auto_out_b_bits_address; // @[BaseTile.scala 190:42]
  wire [7:0] tlMasterXbar_auto_out_b_bits_mask; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_b_bits_corrupt; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_c_ready; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_c_valid; // @[BaseTile.scala 190:42]
  wire [2:0] tlMasterXbar_auto_out_c_bits_opcode; // @[BaseTile.scala 190:42]
  wire [2:0] tlMasterXbar_auto_out_c_bits_param; // @[BaseTile.scala 190:42]
  wire [3:0] tlMasterXbar_auto_out_c_bits_size; // @[BaseTile.scala 190:42]
  wire [1:0] tlMasterXbar_auto_out_c_bits_source; // @[BaseTile.scala 190:42]
  wire [31:0] tlMasterXbar_auto_out_c_bits_address; // @[BaseTile.scala 190:42]
  wire [63:0] tlMasterXbar_auto_out_c_bits_data; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_d_ready; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_d_valid; // @[BaseTile.scala 190:42]
  wire [2:0] tlMasterXbar_auto_out_d_bits_opcode; // @[BaseTile.scala 190:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_param; // @[BaseTile.scala 190:42]
  wire [3:0] tlMasterXbar_auto_out_d_bits_size; // @[BaseTile.scala 190:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_source; // @[BaseTile.scala 190:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_sink; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_d_bits_denied; // @[BaseTile.scala 190:42]
  wire [63:0] tlMasterXbar_auto_out_d_bits_data; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_d_bits_corrupt; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_e_ready; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_auto_out_e_valid; // @[BaseTile.scala 190:42]
  wire [1:0] tlMasterXbar_auto_out_e_bits_sink; // @[BaseTile.scala 190:42]
  wire [29:0] tlMasterXbar_io_covSum; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_metaAssert; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_metaReset; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_TLMonitor_halt; // @[BaseTile.scala 190:42]
  wire  tlMasterXbar_TLMonitor_1_halt; // @[BaseTile.scala 190:42]
  wire  intXbar_auto_int_in_3_0; // @[BaseTile.scala 192:37]
  wire  intXbar_auto_int_in_2_0; // @[BaseTile.scala 192:37]
  wire  intXbar_auto_int_in_1_0; // @[BaseTile.scala 192:37]
  wire  intXbar_auto_int_in_1_1; // @[BaseTile.scala 192:37]
  wire  intXbar_auto_int_in_0_0; // @[BaseTile.scala 192:37]
  wire  intXbar_auto_int_out_0; // @[BaseTile.scala 192:37]
  wire  intXbar_auto_int_out_1; // @[BaseTile.scala 192:37]
  wire  intXbar_auto_int_out_2; // @[BaseTile.scala 192:37]
  wire  intXbar_auto_int_out_3; // @[BaseTile.scala 192:37]
  wire  intXbar_auto_int_out_4; // @[BaseTile.scala 192:37]
  wire [29:0] intXbar_io_covSum; // @[BaseTile.scala 192:37]
  wire  intXbar_metaAssert; // @[BaseTile.scala 192:37]
  wire  hartIdNode_auto_in; // @[BundleBridge.scala 169:31]
  wire  hartIdNode_auto_out_0; // @[BundleBridge.scala 169:31]
  wire [29:0] hartIdNode_io_covSum; // @[BundleBridge.scala 169:31]
  wire  hartIdNode_metaAssert; // @[BundleBridge.scala 169:31]
  wire [31:0] resetVectorNode_auto_in; // @[BundleBridge.scala 169:31]
  wire [31:0] resetVectorNode_auto_out_1; // @[BundleBridge.scala 169:31]
  wire [29:0] resetVectorNode_io_covSum; // @[BundleBridge.scala 169:31]
  wire  resetVectorNode_metaAssert; // @[BundleBridge.scala 169:31]
  wire  dcache_gated_clock; // @[HellaCache.scala 254:43]
  wire  dcache_reset; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_a_ready; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_a_valid; // @[HellaCache.scala 254:43]
  wire [2:0] dcache_auto_out_a_bits_opcode; // @[HellaCache.scala 254:43]
  wire [2:0] dcache_auto_out_a_bits_param; // @[HellaCache.scala 254:43]
  wire [3:0] dcache_auto_out_a_bits_size; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_a_bits_source; // @[HellaCache.scala 254:43]
  wire [31:0] dcache_auto_out_a_bits_address; // @[HellaCache.scala 254:43]
  wire [7:0] dcache_auto_out_a_bits_mask; // @[HellaCache.scala 254:43]
  wire [63:0] dcache_auto_out_a_bits_data; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_b_ready; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_b_valid; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_auto_out_b_bits_param; // @[HellaCache.scala 254:43]
  wire [3:0] dcache_auto_out_b_bits_size; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_b_bits_source; // @[HellaCache.scala 254:43]
  wire [31:0] dcache_auto_out_b_bits_address; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_c_ready; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_c_valid; // @[HellaCache.scala 254:43]
  wire [2:0] dcache_auto_out_c_bits_opcode; // @[HellaCache.scala 254:43]
  wire [2:0] dcache_auto_out_c_bits_param; // @[HellaCache.scala 254:43]
  wire [3:0] dcache_auto_out_c_bits_size; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_c_bits_source; // @[HellaCache.scala 254:43]
  wire [31:0] dcache_auto_out_c_bits_address; // @[HellaCache.scala 254:43]
  wire [63:0] dcache_auto_out_c_bits_data; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_d_ready; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_d_valid; // @[HellaCache.scala 254:43]
  wire [2:0] dcache_auto_out_d_bits_opcode; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_auto_out_d_bits_param; // @[HellaCache.scala 254:43]
  wire [3:0] dcache_auto_out_d_bits_size; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_d_bits_source; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_auto_out_d_bits_sink; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_d_bits_denied; // @[HellaCache.scala 254:43]
  wire [63:0] dcache_auto_out_d_bits_data; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_e_ready; // @[HellaCache.scala 254:43]
  wire  dcache_auto_out_e_valid; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_auto_out_e_bits_sink; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_req_ready; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_req_valid; // @[HellaCache.scala 254:43]
  wire [39:0] dcache_io_cpu_req_bits_addr; // @[HellaCache.scala 254:43]
  wire [6:0] dcache_io_cpu_req_bits_tag; // @[HellaCache.scala 254:43]
  wire [4:0] dcache_io_cpu_req_bits_cmd; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_io_cpu_req_bits_size; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_req_bits_signed; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_req_bits_phys; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_s1_kill; // @[HellaCache.scala 254:43]
  wire [63:0] dcache_io_cpu_s1_data_data; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_s2_nack; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_resp_valid; // @[HellaCache.scala 254:43]
  wire [6:0] dcache_io_cpu_resp_bits_tag; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_io_cpu_resp_bits_size; // @[HellaCache.scala 254:43]
  wire [63:0] dcache_io_cpu_resp_bits_data; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_resp_bits_replay; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_resp_bits_has_data; // @[HellaCache.scala 254:43]
  wire [63:0] dcache_io_cpu_resp_bits_data_word_bypass; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_replay_next; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_s2_xcpt_ma_ld; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_s2_xcpt_ma_st; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_s2_xcpt_pf_ld; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_s2_xcpt_pf_st; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_s2_xcpt_ae_ld; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_s2_xcpt_ae_st; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_ordered; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_perf_release; // @[HellaCache.scala 254:43]
  wire  dcache_io_cpu_perf_grant; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_req_ready; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_req_valid; // @[HellaCache.scala 254:43]
  wire [26:0] dcache_io_ptw_req_bits_bits_addr; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_resp_valid; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_resp_bits_ae; // @[HellaCache.scala 254:43]
  wire [53:0] dcache_io_ptw_resp_bits_pte_ppn; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_resp_bits_pte_d; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_resp_bits_pte_a; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_resp_bits_pte_g; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_resp_bits_pte_u; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_resp_bits_pte_x; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_resp_bits_pte_w; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_resp_bits_pte_r; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_resp_bits_pte_v; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_io_ptw_resp_bits_level; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_resp_bits_homogeneous; // @[HellaCache.scala 254:43]
  wire [3:0] dcache_io_ptw_ptbr_mode; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_status_debug; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_io_ptw_status_dprv; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_status_mxr; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_status_sum; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_0_cfg_l; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_io_ptw_pmp_0_cfg_a; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_0_cfg_x; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_0_cfg_w; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_0_cfg_r; // @[HellaCache.scala 254:43]
  wire [29:0] dcache_io_ptw_pmp_0_addr; // @[HellaCache.scala 254:43]
  wire [31:0] dcache_io_ptw_pmp_0_mask; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_1_cfg_l; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_io_ptw_pmp_1_cfg_a; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_1_cfg_x; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_1_cfg_w; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_1_cfg_r; // @[HellaCache.scala 254:43]
  wire [29:0] dcache_io_ptw_pmp_1_addr; // @[HellaCache.scala 254:43]
  wire [31:0] dcache_io_ptw_pmp_1_mask; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_2_cfg_l; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_io_ptw_pmp_2_cfg_a; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_2_cfg_x; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_2_cfg_w; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_2_cfg_r; // @[HellaCache.scala 254:43]
  wire [29:0] dcache_io_ptw_pmp_2_addr; // @[HellaCache.scala 254:43]
  wire [31:0] dcache_io_ptw_pmp_2_mask; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_3_cfg_l; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_io_ptw_pmp_3_cfg_a; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_3_cfg_x; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_3_cfg_w; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_3_cfg_r; // @[HellaCache.scala 254:43]
  wire [29:0] dcache_io_ptw_pmp_3_addr; // @[HellaCache.scala 254:43]
  wire [31:0] dcache_io_ptw_pmp_3_mask; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_4_cfg_l; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_io_ptw_pmp_4_cfg_a; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_4_cfg_x; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_4_cfg_w; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_4_cfg_r; // @[HellaCache.scala 254:43]
  wire [29:0] dcache_io_ptw_pmp_4_addr; // @[HellaCache.scala 254:43]
  wire [31:0] dcache_io_ptw_pmp_4_mask; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_5_cfg_l; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_io_ptw_pmp_5_cfg_a; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_5_cfg_x; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_5_cfg_w; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_5_cfg_r; // @[HellaCache.scala 254:43]
  wire [29:0] dcache_io_ptw_pmp_5_addr; // @[HellaCache.scala 254:43]
  wire [31:0] dcache_io_ptw_pmp_5_mask; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_6_cfg_l; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_io_ptw_pmp_6_cfg_a; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_6_cfg_x; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_6_cfg_w; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_6_cfg_r; // @[HellaCache.scala 254:43]
  wire [29:0] dcache_io_ptw_pmp_6_addr; // @[HellaCache.scala 254:43]
  wire [31:0] dcache_io_ptw_pmp_6_mask; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_7_cfg_l; // @[HellaCache.scala 254:43]
  wire [1:0] dcache_io_ptw_pmp_7_cfg_a; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_7_cfg_x; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_7_cfg_w; // @[HellaCache.scala 254:43]
  wire  dcache_io_ptw_pmp_7_cfg_r; // @[HellaCache.scala 254:43]
  wire [29:0] dcache_io_ptw_pmp_7_addr; // @[HellaCache.scala 254:43]
  wire [31:0] dcache_io_ptw_pmp_7_mask; // @[HellaCache.scala 254:43]
  wire [29:0] dcache_io_covSum; // @[HellaCache.scala 254:43]
  wire  dcache_metaAssert; // @[HellaCache.scala 254:43]
  wire  dcache_metaReset; // @[HellaCache.scala 254:43]
  wire  dcache_MaxPeriodFibonacciLFSR_halt; // @[HellaCache.scala 254:43]
  wire  dcache_pma_checker_halt; // @[HellaCache.scala 254:43]
  wire  dcache_tlb_halt; // @[HellaCache.scala 254:43]
  wire  dcache_data_halt; // @[HellaCache.scala 254:43]
  wire  frontend_gated_clock; // @[Frontend.scala 352:28]
  wire  frontend_reset; // @[Frontend.scala 352:28]
  wire  frontend_auto_icache_master_out_a_ready; // @[Frontend.scala 352:28]
  wire  frontend_auto_icache_master_out_a_valid; // @[Frontend.scala 352:28]
  wire [31:0] frontend_auto_icache_master_out_a_bits_address; // @[Frontend.scala 352:28]
  wire  frontend_auto_icache_master_out_d_valid; // @[Frontend.scala 352:28]
  wire [2:0] frontend_auto_icache_master_out_d_bits_opcode; // @[Frontend.scala 352:28]
  wire [3:0] frontend_auto_icache_master_out_d_bits_size; // @[Frontend.scala 352:28]
  wire [63:0] frontend_auto_icache_master_out_d_bits_data; // @[Frontend.scala 352:28]
  wire  frontend_auto_icache_master_out_d_bits_corrupt; // @[Frontend.scala 352:28]
  wire [31:0] frontend_auto_reset_vector_sink_in; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_might_request; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_req_valid; // @[Frontend.scala 352:28]
  wire [39:0] frontend_io_cpu_req_bits_pc; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_req_bits_speculative; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_sfence_valid; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_sfence_bits_rs1; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_sfence_bits_rs2; // @[Frontend.scala 352:28]
  wire [38:0] frontend_io_cpu_sfence_bits_addr; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_resp_ready; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_resp_valid; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_resp_bits_btb_taken; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_resp_bits_btb_bridx; // @[Frontend.scala 352:28]
  wire [4:0] frontend_io_cpu_resp_bits_btb_entry; // @[Frontend.scala 352:28]
  wire [7:0] frontend_io_cpu_resp_bits_btb_bht_history; // @[Frontend.scala 352:28]
  wire [39:0] frontend_io_cpu_resp_bits_pc; // @[Frontend.scala 352:28]
  wire [31:0] frontend_io_cpu_resp_bits_data; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_resp_bits_xcpt_pf_inst; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_resp_bits_xcpt_ae_inst; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_resp_bits_replay; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_btb_update_valid; // @[Frontend.scala 352:28]
  wire [4:0] frontend_io_cpu_btb_update_bits_prediction_entry; // @[Frontend.scala 352:28]
  wire [38:0] frontend_io_cpu_btb_update_bits_pc; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_btb_update_bits_isValid; // @[Frontend.scala 352:28]
  wire [38:0] frontend_io_cpu_btb_update_bits_br_pc; // @[Frontend.scala 352:28]
  wire [1:0] frontend_io_cpu_btb_update_bits_cfiType; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_bht_update_valid; // @[Frontend.scala 352:28]
  wire [7:0] frontend_io_cpu_bht_update_bits_prediction_history; // @[Frontend.scala 352:28]
  wire [38:0] frontend_io_cpu_bht_update_bits_pc; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_bht_update_bits_branch; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_bht_update_bits_taken; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_bht_update_bits_mispredict; // @[Frontend.scala 352:28]
  wire  frontend_io_cpu_flush_icache; // @[Frontend.scala 352:28]
  wire [39:0] frontend_io_cpu_npc; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_req_ready; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_req_valid; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_req_bits_valid; // @[Frontend.scala 352:28]
  wire [26:0] frontend_io_ptw_req_bits_bits_addr; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_resp_valid; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_resp_bits_ae; // @[Frontend.scala 352:28]
  wire [53:0] frontend_io_ptw_resp_bits_pte_ppn; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_resp_bits_pte_d; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_resp_bits_pte_a; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_resp_bits_pte_g; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_resp_bits_pte_u; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_resp_bits_pte_x; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_resp_bits_pte_w; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_resp_bits_pte_r; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_resp_bits_pte_v; // @[Frontend.scala 352:28]
  wire [1:0] frontend_io_ptw_resp_bits_level; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_resp_bits_homogeneous; // @[Frontend.scala 352:28]
  wire [3:0] frontend_io_ptw_ptbr_mode; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_status_debug; // @[Frontend.scala 352:28]
  wire [1:0] frontend_io_ptw_status_prv; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_0_cfg_l; // @[Frontend.scala 352:28]
  wire [1:0] frontend_io_ptw_pmp_0_cfg_a; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_0_cfg_x; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_0_cfg_w; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_0_cfg_r; // @[Frontend.scala 352:28]
  wire [29:0] frontend_io_ptw_pmp_0_addr; // @[Frontend.scala 352:28]
  wire [31:0] frontend_io_ptw_pmp_0_mask; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_1_cfg_l; // @[Frontend.scala 352:28]
  wire [1:0] frontend_io_ptw_pmp_1_cfg_a; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_1_cfg_x; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_1_cfg_w; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_1_cfg_r; // @[Frontend.scala 352:28]
  wire [29:0] frontend_io_ptw_pmp_1_addr; // @[Frontend.scala 352:28]
  wire [31:0] frontend_io_ptw_pmp_1_mask; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_2_cfg_l; // @[Frontend.scala 352:28]
  wire [1:0] frontend_io_ptw_pmp_2_cfg_a; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_2_cfg_x; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_2_cfg_w; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_2_cfg_r; // @[Frontend.scala 352:28]
  wire [29:0] frontend_io_ptw_pmp_2_addr; // @[Frontend.scala 352:28]
  wire [31:0] frontend_io_ptw_pmp_2_mask; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_3_cfg_l; // @[Frontend.scala 352:28]
  wire [1:0] frontend_io_ptw_pmp_3_cfg_a; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_3_cfg_x; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_3_cfg_w; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_3_cfg_r; // @[Frontend.scala 352:28]
  wire [29:0] frontend_io_ptw_pmp_3_addr; // @[Frontend.scala 352:28]
  wire [31:0] frontend_io_ptw_pmp_3_mask; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_4_cfg_l; // @[Frontend.scala 352:28]
  wire [1:0] frontend_io_ptw_pmp_4_cfg_a; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_4_cfg_x; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_4_cfg_w; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_4_cfg_r; // @[Frontend.scala 352:28]
  wire [29:0] frontend_io_ptw_pmp_4_addr; // @[Frontend.scala 352:28]
  wire [31:0] frontend_io_ptw_pmp_4_mask; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_5_cfg_l; // @[Frontend.scala 352:28]
  wire [1:0] frontend_io_ptw_pmp_5_cfg_a; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_5_cfg_x; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_5_cfg_w; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_5_cfg_r; // @[Frontend.scala 352:28]
  wire [29:0] frontend_io_ptw_pmp_5_addr; // @[Frontend.scala 352:28]
  wire [31:0] frontend_io_ptw_pmp_5_mask; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_6_cfg_l; // @[Frontend.scala 352:28]
  wire [1:0] frontend_io_ptw_pmp_6_cfg_a; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_6_cfg_x; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_6_cfg_w; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_6_cfg_r; // @[Frontend.scala 352:28]
  wire [29:0] frontend_io_ptw_pmp_6_addr; // @[Frontend.scala 352:28]
  wire [31:0] frontend_io_ptw_pmp_6_mask; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_7_cfg_l; // @[Frontend.scala 352:28]
  wire [1:0] frontend_io_ptw_pmp_7_cfg_a; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_7_cfg_x; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_7_cfg_w; // @[Frontend.scala 352:28]
  wire  frontend_io_ptw_pmp_7_cfg_r; // @[Frontend.scala 352:28]
  wire [29:0] frontend_io_ptw_pmp_7_addr; // @[Frontend.scala 352:28]
  wire [31:0] frontend_io_ptw_pmp_7_mask; // @[Frontend.scala 352:28]
  wire [63:0] frontend_io_ptw_customCSRs_csrs_0_value; // @[Frontend.scala 352:28]
  wire [29:0] frontend_io_covSum; // @[Frontend.scala 352:28]
  wire  frontend_metaAssert; // @[Frontend.scala 352:28]
  wire  frontend_metaReset; // @[Frontend.scala 352:28]
  wire  frontend_icache_halt; // @[Frontend.scala 352:28]
  wire  frontend_fq_halt; // @[Frontend.scala 352:28]
  wire  frontend_tlb_halt; // @[Frontend.scala 352:28]
  wire  frontend_btb_halt; // @[Frontend.scala 352:28]
  wire  buffer_clock; // @[Buffer.scala 69:28]
  wire  buffer_reset; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_a_bits_address; // @[Buffer.scala 69:28]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_a_bits_data; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_a_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_b_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_b_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_b_bits_opcode; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_b_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_in_b_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_b_bits_source; // @[Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_b_bits_address; // @[Buffer.scala 69:28]
  wire [7:0] buffer_auto_in_b_bits_mask; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_b_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_c_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_c_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_c_bits_opcode; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_c_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_in_c_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_c_bits_source; // @[Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_c_bits_address; // @[Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_c_bits_data; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_sink; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_e_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_e_valid; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_e_bits_sink; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_a_bits_address; // @[Buffer.scala 69:28]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_a_bits_data; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_a_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_b_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_b_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_b_bits_opcode; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_b_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_out_b_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_b_bits_source; // @[Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_b_bits_address; // @[Buffer.scala 69:28]
  wire [7:0] buffer_auto_out_b_bits_mask; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_b_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_c_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_c_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_c_bits_opcode; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_c_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_out_c_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_c_bits_source; // @[Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_c_bits_address; // @[Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_c_bits_data; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_c_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_sink; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_d_bits_denied; // @[Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_d_bits_data; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_d_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_e_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_e_valid; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_e_bits_sink; // @[Buffer.scala 69:28]
  wire [29:0] buffer_io_covSum; // @[Buffer.scala 69:28]
  wire  buffer_metaAssert; // @[Buffer.scala 69:28]
  wire  buffer_metaReset; // @[Buffer.scala 69:28]
  wire  buffer_Queue_3_halt; // @[Buffer.scala 69:28]
  wire  buffer_Queue_halt; // @[Buffer.scala 69:28]
  wire  buffer_TLMonitor_halt; // @[Buffer.scala 69:28]
  wire  buffer_Queue_2_halt; // @[Buffer.scala 69:28]
  wire  buffer_Queue_4_halt; // @[Buffer.scala 69:28]
  wire  buffer_Queue_1_halt; // @[Buffer.scala 69:28]
  wire  intsink_clock; // @[Crossing.scala 74:29]
  wire  intsink_auto_in_sync_0; // @[Crossing.scala 74:29]
  wire  intsink_auto_out_0; // @[Crossing.scala 74:29]
  wire [29:0] intsink_io_covSum; // @[Crossing.scala 74:29]
  wire  intsink_metaAssert; // @[Crossing.scala 74:29]
  wire  intsink_metaReset; // @[Crossing.scala 74:29]
  wire  intsink_SynchronizerShiftReg_w1_d3_halt; // @[Crossing.scala 74:29]
  wire  intsink_1_auto_in_sync_0; // @[Crossing.scala 94:29]
  wire  intsink_1_auto_in_sync_1; // @[Crossing.scala 94:29]
  wire  intsink_1_auto_out_0; // @[Crossing.scala 94:29]
  wire  intsink_1_auto_out_1; // @[Crossing.scala 94:29]
  wire [29:0] intsink_1_io_covSum; // @[Crossing.scala 94:29]
  wire  intsink_1_metaAssert; // @[Crossing.scala 94:29]
  wire  intsink_2_auto_in_sync_0; // @[Crossing.scala 94:29]
  wire  intsink_2_auto_out_0; // @[Crossing.scala 94:29]
  wire [29:0] intsink_2_io_covSum; // @[Crossing.scala 94:29]
  wire  intsink_2_metaAssert; // @[Crossing.scala 94:29]
  wire  intsink_3_auto_in_sync_0; // @[Crossing.scala 94:29]
  wire  intsink_3_auto_out_0; // @[Crossing.scala 94:29]
  wire [29:0] intsink_3_io_covSum; // @[Crossing.scala 94:29]
  wire  intsink_3_metaAssert; // @[Crossing.scala 94:29]
  wire  fpuOpt_clock; // @[RocketTile.scala 195:62]
  wire  fpuOpt_reset; // @[RocketTile.scala 195:62]
  wire [31:0] fpuOpt_io_inst; // @[RocketTile.scala 195:62]
  wire [63:0] fpuOpt_io_fromint_data; // @[RocketTile.scala 195:62]
  wire [2:0] fpuOpt_io_fcsr_rm; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_fcsr_flags_valid; // @[RocketTile.scala 195:62]
  wire [4:0] fpuOpt_io_fcsr_flags_bits; // @[RocketTile.scala 195:62]
  wire [63:0] fpuOpt_io_store_data; // @[RocketTile.scala 195:62]
  wire [63:0] fpuOpt_io_toint_data; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_dmem_resp_val; // @[RocketTile.scala 195:62]
  wire [2:0] fpuOpt_io_dmem_resp_type; // @[RocketTile.scala 195:62]
  wire [4:0] fpuOpt_io_dmem_resp_tag; // @[RocketTile.scala 195:62]
  wire [63:0] fpuOpt_io_dmem_resp_data; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_valid; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_fcsr_rdy; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_nack_mem; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_illegal_rm; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_killx; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_killm; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_dec_wen; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_dec_ren1; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_dec_ren2; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_dec_ren3; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_sboard_set; // @[RocketTile.scala 195:62]
  wire  fpuOpt_io_sboard_clr; // @[RocketTile.scala 195:62]
  wire [4:0] fpuOpt_io_sboard_clra; // @[RocketTile.scala 195:62]
  wire [29:0] fpuOpt_io_covSum; // @[RocketTile.scala 195:62]
  wire  fpuOpt_metaAssert; // @[RocketTile.scala 195:62]
  wire  fpuOpt_metaReset; // @[RocketTile.scala 195:62]
  wire  fpuOpt_divSqrt_1_halt; // @[RocketTile.scala 195:62]
  wire  fpuOpt_ifpu_halt; // @[RocketTile.scala 195:62]
  wire  fpuOpt_divSqrt_halt; // @[RocketTile.scala 195:62]
  wire  fpuOpt_fpmu_halt; // @[RocketTile.scala 195:62]
  wire  fpuOpt_dfma_halt; // @[RocketTile.scala 195:62]
  wire  fpuOpt_fpiu_halt; // @[RocketTile.scala 195:62]
  wire  fpuOpt_sfma_halt; // @[RocketTile.scala 195:62]
  wire  dcacheArb_clock; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_0_req_ready; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_0_req_valid; // @[HellaCache.scala 264:25]
  wire [39:0] dcacheArb_io_requestor_0_req_bits_addr; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_0_s1_kill; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_0_s2_nack; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_0_resp_valid; // @[HellaCache.scala 264:25]
  wire [63:0] dcacheArb_io_requestor_0_resp_bits_data; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_0_s2_xcpt_ae_ld; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_req_ready; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_req_valid; // @[HellaCache.scala 264:25]
  wire [39:0] dcacheArb_io_requestor_1_req_bits_addr; // @[HellaCache.scala 264:25]
  wire [6:0] dcacheArb_io_requestor_1_req_bits_tag; // @[HellaCache.scala 264:25]
  wire [4:0] dcacheArb_io_requestor_1_req_bits_cmd; // @[HellaCache.scala 264:25]
  wire [1:0] dcacheArb_io_requestor_1_req_bits_size; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_req_bits_signed; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_s1_kill; // @[HellaCache.scala 264:25]
  wire [63:0] dcacheArb_io_requestor_1_s1_data_data; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_s2_nack; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_resp_valid; // @[HellaCache.scala 264:25]
  wire [6:0] dcacheArb_io_requestor_1_resp_bits_tag; // @[HellaCache.scala 264:25]
  wire [1:0] dcacheArb_io_requestor_1_resp_bits_size; // @[HellaCache.scala 264:25]
  wire [63:0] dcacheArb_io_requestor_1_resp_bits_data; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_resp_bits_replay; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_resp_bits_has_data; // @[HellaCache.scala 264:25]
  wire [63:0] dcacheArb_io_requestor_1_resp_bits_data_word_bypass; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_replay_next; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ma_ld; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ma_st; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_pf_ld; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_pf_st; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ae_ld; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ae_st; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_ordered; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_perf_release; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_requestor_1_perf_grant; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_req_ready; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_req_valid; // @[HellaCache.scala 264:25]
  wire [39:0] dcacheArb_io_mem_req_bits_addr; // @[HellaCache.scala 264:25]
  wire [6:0] dcacheArb_io_mem_req_bits_tag; // @[HellaCache.scala 264:25]
  wire [4:0] dcacheArb_io_mem_req_bits_cmd; // @[HellaCache.scala 264:25]
  wire [1:0] dcacheArb_io_mem_req_bits_size; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_req_bits_signed; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_req_bits_phys; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_s1_kill; // @[HellaCache.scala 264:25]
  wire [63:0] dcacheArb_io_mem_s1_data_data; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_s2_nack; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_resp_valid; // @[HellaCache.scala 264:25]
  wire [6:0] dcacheArb_io_mem_resp_bits_tag; // @[HellaCache.scala 264:25]
  wire [1:0] dcacheArb_io_mem_resp_bits_size; // @[HellaCache.scala 264:25]
  wire [63:0] dcacheArb_io_mem_resp_bits_data; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_resp_bits_replay; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_resp_bits_has_data; // @[HellaCache.scala 264:25]
  wire [63:0] dcacheArb_io_mem_resp_bits_data_word_bypass; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_replay_next; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_s2_xcpt_ma_ld; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_s2_xcpt_ma_st; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_s2_xcpt_pf_ld; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_s2_xcpt_pf_st; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_s2_xcpt_ae_ld; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_s2_xcpt_ae_st; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_ordered; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_perf_release; // @[HellaCache.scala 264:25]
  wire  dcacheArb_io_mem_perf_grant; // @[HellaCache.scala 264:25]
  wire [29:0] dcacheArb_io_covSum; // @[HellaCache.scala 264:25]
  wire  dcacheArb_metaAssert; // @[HellaCache.scala 264:25]
  wire  dcacheArb_metaReset; // @[HellaCache.scala 264:25]
  wire  ptw_clock; // @[PTW.scala 395:19]
  wire  ptw_reset; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_req_ready; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_req_valid; // @[PTW.scala 395:19]
  wire [26:0] ptw_io_requestor_0_req_bits_bits_addr; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_resp_valid; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_resp_bits_ae; // @[PTW.scala 395:19]
  wire [53:0] ptw_io_requestor_0_resp_bits_pte_ppn; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_resp_bits_pte_d; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_resp_bits_pte_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_resp_bits_pte_g; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_resp_bits_pte_u; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_resp_bits_pte_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_resp_bits_pte_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_resp_bits_pte_r; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_resp_bits_pte_v; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_0_resp_bits_level; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_resp_bits_homogeneous; // @[PTW.scala 395:19]
  wire [3:0] ptw_io_requestor_0_ptbr_mode; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_status_debug; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_0_status_dprv; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_status_mxr; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_status_sum; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_0_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_0_pmp_0_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_0_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_0_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_0_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_0_pmp_0_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_0_pmp_0_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_1_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_0_pmp_1_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_1_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_1_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_1_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_0_pmp_1_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_0_pmp_1_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_2_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_0_pmp_2_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_2_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_2_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_2_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_0_pmp_2_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_0_pmp_2_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_3_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_0_pmp_3_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_3_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_3_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_3_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_0_pmp_3_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_0_pmp_3_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_4_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_0_pmp_4_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_4_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_4_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_4_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_0_pmp_4_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_0_pmp_4_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_5_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_0_pmp_5_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_5_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_5_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_5_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_0_pmp_5_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_0_pmp_5_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_6_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_0_pmp_6_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_6_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_6_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_6_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_0_pmp_6_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_0_pmp_6_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_7_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_0_pmp_7_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_7_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_7_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_0_pmp_7_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_0_pmp_7_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_0_pmp_7_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_req_ready; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_req_valid; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_req_bits_valid; // @[PTW.scala 395:19]
  wire [26:0] ptw_io_requestor_1_req_bits_bits_addr; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_resp_valid; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_resp_bits_ae; // @[PTW.scala 395:19]
  wire [53:0] ptw_io_requestor_1_resp_bits_pte_ppn; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_resp_bits_pte_d; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_resp_bits_pte_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_resp_bits_pte_g; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_resp_bits_pte_u; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_resp_bits_pte_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_resp_bits_pte_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_resp_bits_pte_r; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_resp_bits_pte_v; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_1_resp_bits_level; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_resp_bits_homogeneous; // @[PTW.scala 395:19]
  wire [3:0] ptw_io_requestor_1_ptbr_mode; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_status_debug; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_1_status_prv; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_0_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_1_pmp_0_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_0_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_0_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_0_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_1_pmp_0_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_1_pmp_0_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_1_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_1_pmp_1_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_1_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_1_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_1_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_1_pmp_1_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_1_pmp_1_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_2_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_1_pmp_2_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_2_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_2_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_2_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_1_pmp_2_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_1_pmp_2_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_3_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_1_pmp_3_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_3_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_3_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_3_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_1_pmp_3_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_1_pmp_3_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_4_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_1_pmp_4_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_4_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_4_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_4_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_1_pmp_4_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_1_pmp_4_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_5_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_1_pmp_5_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_5_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_5_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_5_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_1_pmp_5_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_1_pmp_5_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_6_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_1_pmp_6_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_6_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_6_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_6_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_1_pmp_6_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_1_pmp_6_mask; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_7_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_requestor_1_pmp_7_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_7_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_7_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_requestor_1_pmp_7_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_requestor_1_pmp_7_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_requestor_1_pmp_7_mask; // @[PTW.scala 395:19]
  wire [63:0] ptw_io_requestor_1_customCSRs_csrs_0_value; // @[PTW.scala 395:19]
  wire  ptw_io_mem_req_ready; // @[PTW.scala 395:19]
  wire  ptw_io_mem_req_valid; // @[PTW.scala 395:19]
  wire [39:0] ptw_io_mem_req_bits_addr; // @[PTW.scala 395:19]
  wire  ptw_io_mem_s1_kill; // @[PTW.scala 395:19]
  wire  ptw_io_mem_s2_nack; // @[PTW.scala 395:19]
  wire  ptw_io_mem_resp_valid; // @[PTW.scala 395:19]
  wire [63:0] ptw_io_mem_resp_bits_data; // @[PTW.scala 395:19]
  wire  ptw_io_mem_s2_xcpt_ae_ld; // @[PTW.scala 395:19]
  wire [3:0] ptw_io_dpath_ptbr_mode; // @[PTW.scala 395:19]
  wire [43:0] ptw_io_dpath_ptbr_ppn; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_sfence_valid; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_sfence_bits_rs1; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_status_debug; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_dpath_status_dprv; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_dpath_status_prv; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_status_mxr; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_status_sum; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_0_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_dpath_pmp_0_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_0_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_0_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_0_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_dpath_pmp_0_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_dpath_pmp_0_mask; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_1_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_dpath_pmp_1_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_1_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_1_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_1_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_dpath_pmp_1_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_dpath_pmp_1_mask; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_2_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_dpath_pmp_2_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_2_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_2_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_2_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_dpath_pmp_2_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_dpath_pmp_2_mask; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_3_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_dpath_pmp_3_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_3_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_3_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_3_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_dpath_pmp_3_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_dpath_pmp_3_mask; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_4_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_dpath_pmp_4_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_4_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_4_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_4_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_dpath_pmp_4_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_dpath_pmp_4_mask; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_5_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_dpath_pmp_5_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_5_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_5_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_5_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_dpath_pmp_5_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_dpath_pmp_5_mask; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_6_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_dpath_pmp_6_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_6_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_6_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_6_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_dpath_pmp_6_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_dpath_pmp_6_mask; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_7_cfg_l; // @[PTW.scala 395:19]
  wire [1:0] ptw_io_dpath_pmp_7_cfg_a; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_7_cfg_x; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_7_cfg_w; // @[PTW.scala 395:19]
  wire  ptw_io_dpath_pmp_7_cfg_r; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_dpath_pmp_7_addr; // @[PTW.scala 395:19]
  wire [31:0] ptw_io_dpath_pmp_7_mask; // @[PTW.scala 395:19]
  wire [63:0] ptw_io_dpath_customCSRs_csrs_0_value; // @[PTW.scala 395:19]
  wire [29:0] ptw_io_covSum; // @[PTW.scala 395:19]
  wire  ptw_metaAssert; // @[PTW.scala 395:19]
  wire  ptw_metaReset; // @[PTW.scala 395:19]
  wire  core_clock; // @[RocketTile.scala 135:20]
  wire  core_reset; // @[RocketTile.scala 135:20]
  wire  core_io_hartid; // @[RocketTile.scala 135:20]
  wire  core_io_interrupts_debug; // @[RocketTile.scala 135:20]
  wire  core_io_interrupts_mtip; // @[RocketTile.scala 135:20]
  wire  core_io_interrupts_msip; // @[RocketTile.scala 135:20]
  wire  core_io_interrupts_meip; // @[RocketTile.scala 135:20]
  wire  core_io_interrupts_seip; // @[RocketTile.scala 135:20]
  wire  core_io_imem_might_request; // @[RocketTile.scala 135:20]
  wire  core_io_imem_req_valid; // @[RocketTile.scala 135:20]
  wire [39:0] core_io_imem_req_bits_pc; // @[RocketTile.scala 135:20]
  wire  core_io_imem_req_bits_speculative; // @[RocketTile.scala 135:20]
  wire  core_io_imem_sfence_valid; // @[RocketTile.scala 135:20]
  wire  core_io_imem_sfence_bits_rs1; // @[RocketTile.scala 135:20]
  wire  core_io_imem_sfence_bits_rs2; // @[RocketTile.scala 135:20]
  wire [38:0] core_io_imem_sfence_bits_addr; // @[RocketTile.scala 135:20]
  wire  core_io_imem_resp_ready; // @[RocketTile.scala 135:20]
  wire  core_io_imem_resp_valid; // @[RocketTile.scala 135:20]
  wire  core_io_imem_resp_bits_btb_taken; // @[RocketTile.scala 135:20]
  wire  core_io_imem_resp_bits_btb_bridx; // @[RocketTile.scala 135:20]
  wire [4:0] core_io_imem_resp_bits_btb_entry; // @[RocketTile.scala 135:20]
  wire [7:0] core_io_imem_resp_bits_btb_bht_history; // @[RocketTile.scala 135:20]
  wire [39:0] core_io_imem_resp_bits_pc; // @[RocketTile.scala 135:20]
  wire [31:0] core_io_imem_resp_bits_data; // @[RocketTile.scala 135:20]
  wire  core_io_imem_resp_bits_xcpt_pf_inst; // @[RocketTile.scala 135:20]
  wire  core_io_imem_resp_bits_xcpt_ae_inst; // @[RocketTile.scala 135:20]
  wire  core_io_imem_resp_bits_replay; // @[RocketTile.scala 135:20]
  wire  core_io_imem_btb_update_valid; // @[RocketTile.scala 135:20]
  wire [4:0] core_io_imem_btb_update_bits_prediction_entry; // @[RocketTile.scala 135:20]
  wire [38:0] core_io_imem_btb_update_bits_pc; // @[RocketTile.scala 135:20]
  wire  core_io_imem_btb_update_bits_isValid; // @[RocketTile.scala 135:20]
  wire [38:0] core_io_imem_btb_update_bits_br_pc; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_imem_btb_update_bits_cfiType; // @[RocketTile.scala 135:20]
  wire  core_io_imem_bht_update_valid; // @[RocketTile.scala 135:20]
  wire [7:0] core_io_imem_bht_update_bits_prediction_history; // @[RocketTile.scala 135:20]
  wire [38:0] core_io_imem_bht_update_bits_pc; // @[RocketTile.scala 135:20]
  wire  core_io_imem_bht_update_bits_branch; // @[RocketTile.scala 135:20]
  wire  core_io_imem_bht_update_bits_taken; // @[RocketTile.scala 135:20]
  wire  core_io_imem_bht_update_bits_mispredict; // @[RocketTile.scala 135:20]
  wire  core_io_imem_flush_icache; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_req_ready; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_req_valid; // @[RocketTile.scala 135:20]
  wire [39:0] core_io_dmem_req_bits_addr; // @[RocketTile.scala 135:20]
  wire [6:0] core_io_dmem_req_bits_tag; // @[RocketTile.scala 135:20]
  wire [4:0] core_io_dmem_req_bits_cmd; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_dmem_req_bits_size; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_req_bits_signed; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_s1_kill; // @[RocketTile.scala 135:20]
  wire [63:0] core_io_dmem_s1_data_data; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_s2_nack; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_resp_valid; // @[RocketTile.scala 135:20]
  wire [6:0] core_io_dmem_resp_bits_tag; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_dmem_resp_bits_size; // @[RocketTile.scala 135:20]
  wire [63:0] core_io_dmem_resp_bits_data; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_resp_bits_replay; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_resp_bits_has_data; // @[RocketTile.scala 135:20]
  wire [63:0] core_io_dmem_resp_bits_data_word_bypass; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_replay_next; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_s2_xcpt_ma_ld; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_s2_xcpt_ma_st; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_s2_xcpt_pf_ld; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_s2_xcpt_pf_st; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_s2_xcpt_ae_ld; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_s2_xcpt_ae_st; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_ordered; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_perf_release; // @[RocketTile.scala 135:20]
  wire  core_io_dmem_perf_grant; // @[RocketTile.scala 135:20]
  wire [3:0] core_io_ptw_ptbr_mode; // @[RocketTile.scala 135:20]
  wire [43:0] core_io_ptw_ptbr_ppn; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_sfence_valid; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_sfence_bits_rs1; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_status_debug; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_ptw_status_dprv; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_ptw_status_prv; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_status_mxr; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_status_sum; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_0_cfg_l; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_ptw_pmp_0_cfg_a; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_0_cfg_x; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_0_cfg_w; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_0_cfg_r; // @[RocketTile.scala 135:20]
  wire [29:0] core_io_ptw_pmp_0_addr; // @[RocketTile.scala 135:20]
  wire [31:0] core_io_ptw_pmp_0_mask; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_1_cfg_l; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_ptw_pmp_1_cfg_a; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_1_cfg_x; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_1_cfg_w; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_1_cfg_r; // @[RocketTile.scala 135:20]
  wire [29:0] core_io_ptw_pmp_1_addr; // @[RocketTile.scala 135:20]
  wire [31:0] core_io_ptw_pmp_1_mask; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_2_cfg_l; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_ptw_pmp_2_cfg_a; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_2_cfg_x; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_2_cfg_w; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_2_cfg_r; // @[RocketTile.scala 135:20]
  wire [29:0] core_io_ptw_pmp_2_addr; // @[RocketTile.scala 135:20]
  wire [31:0] core_io_ptw_pmp_2_mask; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_3_cfg_l; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_ptw_pmp_3_cfg_a; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_3_cfg_x; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_3_cfg_w; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_3_cfg_r; // @[RocketTile.scala 135:20]
  wire [29:0] core_io_ptw_pmp_3_addr; // @[RocketTile.scala 135:20]
  wire [31:0] core_io_ptw_pmp_3_mask; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_4_cfg_l; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_ptw_pmp_4_cfg_a; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_4_cfg_x; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_4_cfg_w; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_4_cfg_r; // @[RocketTile.scala 135:20]
  wire [29:0] core_io_ptw_pmp_4_addr; // @[RocketTile.scala 135:20]
  wire [31:0] core_io_ptw_pmp_4_mask; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_5_cfg_l; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_ptw_pmp_5_cfg_a; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_5_cfg_x; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_5_cfg_w; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_5_cfg_r; // @[RocketTile.scala 135:20]
  wire [29:0] core_io_ptw_pmp_5_addr; // @[RocketTile.scala 135:20]
  wire [31:0] core_io_ptw_pmp_5_mask; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_6_cfg_l; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_ptw_pmp_6_cfg_a; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_6_cfg_x; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_6_cfg_w; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_6_cfg_r; // @[RocketTile.scala 135:20]
  wire [29:0] core_io_ptw_pmp_6_addr; // @[RocketTile.scala 135:20]
  wire [31:0] core_io_ptw_pmp_6_mask; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_7_cfg_l; // @[RocketTile.scala 135:20]
  wire [1:0] core_io_ptw_pmp_7_cfg_a; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_7_cfg_x; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_7_cfg_w; // @[RocketTile.scala 135:20]
  wire  core_io_ptw_pmp_7_cfg_r; // @[RocketTile.scala 135:20]
  wire [29:0] core_io_ptw_pmp_7_addr; // @[RocketTile.scala 135:20]
  wire [31:0] core_io_ptw_pmp_7_mask; // @[RocketTile.scala 135:20]
  wire [63:0] core_io_ptw_customCSRs_csrs_0_value; // @[RocketTile.scala 135:20]
  wire [31:0] core_io_fpu_inst; // @[RocketTile.scala 135:20]
  wire [63:0] core_io_fpu_fromint_data; // @[RocketTile.scala 135:20]
  wire [2:0] core_io_fpu_fcsr_rm; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_fcsr_flags_valid; // @[RocketTile.scala 135:20]
  wire [4:0] core_io_fpu_fcsr_flags_bits; // @[RocketTile.scala 135:20]
  wire [63:0] core_io_fpu_store_data; // @[RocketTile.scala 135:20]
  wire [63:0] core_io_fpu_toint_data; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_dmem_resp_val; // @[RocketTile.scala 135:20]
  wire [2:0] core_io_fpu_dmem_resp_type; // @[RocketTile.scala 135:20]
  wire [4:0] core_io_fpu_dmem_resp_tag; // @[RocketTile.scala 135:20]
  wire [63:0] core_io_fpu_dmem_resp_data; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_valid; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_fcsr_rdy; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_nack_mem; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_illegal_rm; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_killx; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_killm; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_dec_wen; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_dec_ren1; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_dec_ren2; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_dec_ren3; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_sboard_set; // @[RocketTile.scala 135:20]
  wire  core_io_fpu_sboard_clr; // @[RocketTile.scala 135:20]
  wire [4:0] core_io_fpu_sboard_clra; // @[RocketTile.scala 135:20]
  wire  core_io_wfi; // @[RocketTile.scala 135:20]
  wire [29:0] core_io_covSum; // @[RocketTile.scala 135:20]
  wire  core_metaAssert; // @[RocketTile.scala 135:20]
  wire  core_metaReset; // @[RocketTile.scala 135:20]
  wire  core_csr_halt; // @[RocketTile.scala 135:20]
  wire  core_div_halt; // @[RocketTile.scala 135:20]
  wire  core_ibuf_halt; // @[RocketTile.scala 135:20]
  reg  _T_33; // @[Interrupts.scala 119:36]
  reg [31:0] _RAND_0;
  wire [29:0] RocketTile_covSum;
  wire [29:0] ptw_sum;
  wire [29:0] resetVectorNode_sum;
  wire [29:0] dcacheArb_sum;
  wire [29:0] tlMasterXbar_sum;
  wire [29:0] dcache_sum;
  wire [29:0] intsink_3_sum;
  wire [29:0] intsink_1_sum;
  wire [29:0] buffer_sum;
  wire [29:0] core_sum;
  wire [29:0] fpuOpt_sum;
  wire [29:0] intXbar_sum;
  wire [29:0] frontend_sum;
  wire [29:0] hartIdNode_sum;
  wire [29:0] intsink_sum;
  wire [29:0] intsink_2_sum;
  wire  ptw_metaAssert_wire;
  wire  intsink_2_metaAssert_wire;
  wire  hartIdNode_metaAssert_wire;
  wire  intsink_metaAssert_wire;
  wire  fpuOpt_metaAssert_wire;
  wire  resetVectorNode_metaAssert_wire;
  wire  frontend_metaAssert_wire;
  wire  dcacheArb_metaAssert_wire;
  wire  buffer_metaAssert_wire;
  wire  intsink_1_metaAssert_wire;
  wire  intXbar_metaAssert_wire;
  wire  core_metaAssert_wire;
  wire  tlMasterXbar_metaAssert_wire;
  wire  intsink_3_metaAssert_wire;
  wire  dcache_metaAssert_wire;
  wire  RocketTile_or8;
  wire  RocketTile_or3;
  wire  RocketTile_or9;
  wire  RocketTile_or10;
  wire  RocketTile_or4;
  wire  RocketTile_or1;
  wire  RocketTile_or11;
  wire  RocketTile_or12;
  wire  RocketTile_or5;
  wire  RocketTile_or13;
  wire  RocketTile_or14;
  wire  RocketTile_or6;
  wire  RocketTile_or2;
  wire  RocketTile_or0;
  reg  RocketTile_metaAssert;
  reg [31:0] _RAND_1;
  TLXbar_7 tlMasterXbar ( // @[BaseTile.scala 190:42]
    .clock(tlMasterXbar_clock),
    .reset(tlMasterXbar_reset),
    .auto_in_1_a_ready(tlMasterXbar_auto_in_1_a_ready),
    .auto_in_1_a_valid(tlMasterXbar_auto_in_1_a_valid),
    .auto_in_1_a_bits_address(tlMasterXbar_auto_in_1_a_bits_address),
    .auto_in_1_d_valid(tlMasterXbar_auto_in_1_d_valid),
    .auto_in_1_d_bits_opcode(tlMasterXbar_auto_in_1_d_bits_opcode),
    .auto_in_1_d_bits_size(tlMasterXbar_auto_in_1_d_bits_size),
    .auto_in_1_d_bits_data(tlMasterXbar_auto_in_1_d_bits_data),
    .auto_in_1_d_bits_corrupt(tlMasterXbar_auto_in_1_d_bits_corrupt),
    .auto_in_0_a_ready(tlMasterXbar_auto_in_0_a_ready),
    .auto_in_0_a_valid(tlMasterXbar_auto_in_0_a_valid),
    .auto_in_0_a_bits_opcode(tlMasterXbar_auto_in_0_a_bits_opcode),
    .auto_in_0_a_bits_param(tlMasterXbar_auto_in_0_a_bits_param),
    .auto_in_0_a_bits_size(tlMasterXbar_auto_in_0_a_bits_size),
    .auto_in_0_a_bits_source(tlMasterXbar_auto_in_0_a_bits_source),
    .auto_in_0_a_bits_address(tlMasterXbar_auto_in_0_a_bits_address),
    .auto_in_0_a_bits_mask(tlMasterXbar_auto_in_0_a_bits_mask),
    .auto_in_0_a_bits_data(tlMasterXbar_auto_in_0_a_bits_data),
    .auto_in_0_b_ready(tlMasterXbar_auto_in_0_b_ready),
    .auto_in_0_b_valid(tlMasterXbar_auto_in_0_b_valid),
    .auto_in_0_b_bits_param(tlMasterXbar_auto_in_0_b_bits_param),
    .auto_in_0_b_bits_size(tlMasterXbar_auto_in_0_b_bits_size),
    .auto_in_0_b_bits_source(tlMasterXbar_auto_in_0_b_bits_source),
    .auto_in_0_b_bits_address(tlMasterXbar_auto_in_0_b_bits_address),
    .auto_in_0_c_ready(tlMasterXbar_auto_in_0_c_ready),
    .auto_in_0_c_valid(tlMasterXbar_auto_in_0_c_valid),
    .auto_in_0_c_bits_opcode(tlMasterXbar_auto_in_0_c_bits_opcode),
    .auto_in_0_c_bits_param(tlMasterXbar_auto_in_0_c_bits_param),
    .auto_in_0_c_bits_size(tlMasterXbar_auto_in_0_c_bits_size),
    .auto_in_0_c_bits_source(tlMasterXbar_auto_in_0_c_bits_source),
    .auto_in_0_c_bits_address(tlMasterXbar_auto_in_0_c_bits_address),
    .auto_in_0_c_bits_data(tlMasterXbar_auto_in_0_c_bits_data),
    .auto_in_0_d_ready(tlMasterXbar_auto_in_0_d_ready),
    .auto_in_0_d_valid(tlMasterXbar_auto_in_0_d_valid),
    .auto_in_0_d_bits_opcode(tlMasterXbar_auto_in_0_d_bits_opcode),
    .auto_in_0_d_bits_param(tlMasterXbar_auto_in_0_d_bits_param),
    .auto_in_0_d_bits_size(tlMasterXbar_auto_in_0_d_bits_size),
    .auto_in_0_d_bits_source(tlMasterXbar_auto_in_0_d_bits_source),
    .auto_in_0_d_bits_sink(tlMasterXbar_auto_in_0_d_bits_sink),
    .auto_in_0_d_bits_denied(tlMasterXbar_auto_in_0_d_bits_denied),
    .auto_in_0_d_bits_data(tlMasterXbar_auto_in_0_d_bits_data),
    .auto_in_0_e_ready(tlMasterXbar_auto_in_0_e_ready),
    .auto_in_0_e_valid(tlMasterXbar_auto_in_0_e_valid),
    .auto_in_0_e_bits_sink(tlMasterXbar_auto_in_0_e_bits_sink),
    .auto_out_a_ready(tlMasterXbar_auto_out_a_ready),
    .auto_out_a_valid(tlMasterXbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(tlMasterXbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(tlMasterXbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(tlMasterXbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(tlMasterXbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(tlMasterXbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(tlMasterXbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(tlMasterXbar_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(tlMasterXbar_auto_out_a_bits_corrupt),
    .auto_out_b_ready(tlMasterXbar_auto_out_b_ready),
    .auto_out_b_valid(tlMasterXbar_auto_out_b_valid),
    .auto_out_b_bits_opcode(tlMasterXbar_auto_out_b_bits_opcode),
    .auto_out_b_bits_param(tlMasterXbar_auto_out_b_bits_param),
    .auto_out_b_bits_size(tlMasterXbar_auto_out_b_bits_size),
    .auto_out_b_bits_source(tlMasterXbar_auto_out_b_bits_source),
    .auto_out_b_bits_address(tlMasterXbar_auto_out_b_bits_address),
    .auto_out_b_bits_mask(tlMasterXbar_auto_out_b_bits_mask),
    .auto_out_b_bits_corrupt(tlMasterXbar_auto_out_b_bits_corrupt),
    .auto_out_c_ready(tlMasterXbar_auto_out_c_ready),
    .auto_out_c_valid(tlMasterXbar_auto_out_c_valid),
    .auto_out_c_bits_opcode(tlMasterXbar_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(tlMasterXbar_auto_out_c_bits_param),
    .auto_out_c_bits_size(tlMasterXbar_auto_out_c_bits_size),
    .auto_out_c_bits_source(tlMasterXbar_auto_out_c_bits_source),
    .auto_out_c_bits_address(tlMasterXbar_auto_out_c_bits_address),
    .auto_out_c_bits_data(tlMasterXbar_auto_out_c_bits_data),
    .auto_out_d_ready(tlMasterXbar_auto_out_d_ready),
    .auto_out_d_valid(tlMasterXbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(tlMasterXbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(tlMasterXbar_auto_out_d_bits_param),
    .auto_out_d_bits_size(tlMasterXbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(tlMasterXbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(tlMasterXbar_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(tlMasterXbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(tlMasterXbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(tlMasterXbar_auto_out_d_bits_corrupt),
    .auto_out_e_ready(tlMasterXbar_auto_out_e_ready),
    .auto_out_e_valid(tlMasterXbar_auto_out_e_valid),
    .auto_out_e_bits_sink(tlMasterXbar_auto_out_e_bits_sink),
    .io_covSum(tlMasterXbar_io_covSum),
    .metaAssert(tlMasterXbar_metaAssert),
    .metaReset(tlMasterXbar_metaReset),
    .TLMonitor_halt(tlMasterXbar_TLMonitor_halt),
    .TLMonitor_1_halt(tlMasterXbar_TLMonitor_1_halt)
  );
  IntXbar_1 intXbar ( // @[BaseTile.scala 192:37]
    .auto_int_in_3_0(intXbar_auto_int_in_3_0),
    .auto_int_in_2_0(intXbar_auto_int_in_2_0),
    .auto_int_in_1_0(intXbar_auto_int_in_1_0),
    .auto_int_in_1_1(intXbar_auto_int_in_1_1),
    .auto_int_in_0_0(intXbar_auto_int_in_0_0),
    .auto_int_out_0(intXbar_auto_int_out_0),
    .auto_int_out_1(intXbar_auto_int_out_1),
    .auto_int_out_2(intXbar_auto_int_out_2),
    .auto_int_out_3(intXbar_auto_int_out_3),
    .auto_int_out_4(intXbar_auto_int_out_4),
    .io_covSum(intXbar_io_covSum),
    .metaAssert(intXbar_metaAssert)
  );
  BundleBridgeNexus hartIdNode ( // @[BundleBridge.scala 169:31]
    .auto_in(hartIdNode_auto_in),
    .auto_out_0(hartIdNode_auto_out_0),
    .io_covSum(hartIdNode_io_covSum),
    .metaAssert(hartIdNode_metaAssert)
  );
  BundleBridgeNexus_1 resetVectorNode ( // @[BundleBridge.scala 169:31]
    .auto_in(resetVectorNode_auto_in),
    .auto_out_1(resetVectorNode_auto_out_1),
    .io_covSum(resetVectorNode_io_covSum),
    .metaAssert(resetVectorNode_metaAssert)
  );
  DCache dcache ( // @[HellaCache.scala 254:43]
    .gated_clock(dcache_gated_clock),
    .reset(dcache_reset),
    .auto_out_a_ready(dcache_auto_out_a_ready),
    .auto_out_a_valid(dcache_auto_out_a_valid),
    .auto_out_a_bits_opcode(dcache_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(dcache_auto_out_a_bits_param),
    .auto_out_a_bits_size(dcache_auto_out_a_bits_size),
    .auto_out_a_bits_source(dcache_auto_out_a_bits_source),
    .auto_out_a_bits_address(dcache_auto_out_a_bits_address),
    .auto_out_a_bits_mask(dcache_auto_out_a_bits_mask),
    .auto_out_a_bits_data(dcache_auto_out_a_bits_data),
    .auto_out_b_ready(dcache_auto_out_b_ready),
    .auto_out_b_valid(dcache_auto_out_b_valid),
    .auto_out_b_bits_param(dcache_auto_out_b_bits_param),
    .auto_out_b_bits_size(dcache_auto_out_b_bits_size),
    .auto_out_b_bits_source(dcache_auto_out_b_bits_source),
    .auto_out_b_bits_address(dcache_auto_out_b_bits_address),
    .auto_out_c_ready(dcache_auto_out_c_ready),
    .auto_out_c_valid(dcache_auto_out_c_valid),
    .auto_out_c_bits_opcode(dcache_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(dcache_auto_out_c_bits_param),
    .auto_out_c_bits_size(dcache_auto_out_c_bits_size),
    .auto_out_c_bits_source(dcache_auto_out_c_bits_source),
    .auto_out_c_bits_address(dcache_auto_out_c_bits_address),
    .auto_out_c_bits_data(dcache_auto_out_c_bits_data),
    .auto_out_d_ready(dcache_auto_out_d_ready),
    .auto_out_d_valid(dcache_auto_out_d_valid),
    .auto_out_d_bits_opcode(dcache_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(dcache_auto_out_d_bits_param),
    .auto_out_d_bits_size(dcache_auto_out_d_bits_size),
    .auto_out_d_bits_source(dcache_auto_out_d_bits_source),
    .auto_out_d_bits_sink(dcache_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(dcache_auto_out_d_bits_denied),
    .auto_out_d_bits_data(dcache_auto_out_d_bits_data),
    .auto_out_e_ready(dcache_auto_out_e_ready),
    .auto_out_e_valid(dcache_auto_out_e_valid),
    .auto_out_e_bits_sink(dcache_auto_out_e_bits_sink),
    .io_cpu_req_ready(dcache_io_cpu_req_ready),
    .io_cpu_req_valid(dcache_io_cpu_req_valid),
    .io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr),
    .io_cpu_req_bits_tag(dcache_io_cpu_req_bits_tag),
    .io_cpu_req_bits_cmd(dcache_io_cpu_req_bits_cmd),
    .io_cpu_req_bits_size(dcache_io_cpu_req_bits_size),
    .io_cpu_req_bits_signed(dcache_io_cpu_req_bits_signed),
    .io_cpu_req_bits_phys(dcache_io_cpu_req_bits_phys),
    .io_cpu_s1_kill(dcache_io_cpu_s1_kill),
    .io_cpu_s1_data_data(dcache_io_cpu_s1_data_data),
    .io_cpu_s2_nack(dcache_io_cpu_s2_nack),
    .io_cpu_resp_valid(dcache_io_cpu_resp_valid),
    .io_cpu_resp_bits_tag(dcache_io_cpu_resp_bits_tag),
    .io_cpu_resp_bits_size(dcache_io_cpu_resp_bits_size),
    .io_cpu_resp_bits_data(dcache_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_replay(dcache_io_cpu_resp_bits_replay),
    .io_cpu_resp_bits_has_data(dcache_io_cpu_resp_bits_has_data),
    .io_cpu_resp_bits_data_word_bypass(dcache_io_cpu_resp_bits_data_word_bypass),
    .io_cpu_replay_next(dcache_io_cpu_replay_next),
    .io_cpu_s2_xcpt_ma_ld(dcache_io_cpu_s2_xcpt_ma_ld),
    .io_cpu_s2_xcpt_ma_st(dcache_io_cpu_s2_xcpt_ma_st),
    .io_cpu_s2_xcpt_pf_ld(dcache_io_cpu_s2_xcpt_pf_ld),
    .io_cpu_s2_xcpt_pf_st(dcache_io_cpu_s2_xcpt_pf_st),
    .io_cpu_s2_xcpt_ae_ld(dcache_io_cpu_s2_xcpt_ae_ld),
    .io_cpu_s2_xcpt_ae_st(dcache_io_cpu_s2_xcpt_ae_st),
    .io_cpu_ordered(dcache_io_cpu_ordered),
    .io_cpu_perf_release(dcache_io_cpu_perf_release),
    .io_cpu_perf_grant(dcache_io_cpu_perf_grant),
    .io_ptw_req_ready(dcache_io_ptw_req_ready),
    .io_ptw_req_valid(dcache_io_ptw_req_valid),
    .io_ptw_req_bits_bits_addr(dcache_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(dcache_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(dcache_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(dcache_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(dcache_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(dcache_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(dcache_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(dcache_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(dcache_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(dcache_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(dcache_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(dcache_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(dcache_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(dcache_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(dcache_io_ptw_ptbr_mode),
    .io_ptw_status_debug(dcache_io_ptw_status_debug),
    .io_ptw_status_dprv(dcache_io_ptw_status_dprv),
    .io_ptw_status_mxr(dcache_io_ptw_status_mxr),
    .io_ptw_status_sum(dcache_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(dcache_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(dcache_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(dcache_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(dcache_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(dcache_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(dcache_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(dcache_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(dcache_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(dcache_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(dcache_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(dcache_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(dcache_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(dcache_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(dcache_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(dcache_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(dcache_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(dcache_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(dcache_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(dcache_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(dcache_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(dcache_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(dcache_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(dcache_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(dcache_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(dcache_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(dcache_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(dcache_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(dcache_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(dcache_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(dcache_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(dcache_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(dcache_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(dcache_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(dcache_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(dcache_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(dcache_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(dcache_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(dcache_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(dcache_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(dcache_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(dcache_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(dcache_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(dcache_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(dcache_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(dcache_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(dcache_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(dcache_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(dcache_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(dcache_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(dcache_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(dcache_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(dcache_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(dcache_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(dcache_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(dcache_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(dcache_io_ptw_pmp_7_mask),
    .io_covSum(dcache_io_covSum),
    .metaAssert(dcache_metaAssert),
    .metaReset(dcache_metaReset),
    .MaxPeriodFibonacciLFSR_halt(dcache_MaxPeriodFibonacciLFSR_halt),
    .pma_checker_halt(dcache_pma_checker_halt),
    .tlb_halt(dcache_tlb_halt),
    .data_halt(dcache_data_halt),
    .Checking_DCache_regstate(DCache_regstate),		//Jaewon_DCache_regstate
    .Checking_DCache_covSum(DCache_covSum)			//Jaewon_DCache_regstate
  );
  Frontend frontend ( // @[Frontend.scala 352:28]
	.Checking_Frontend_regstate(Frontend_regstate), 	//Jaewon_regstate
	.Checking_Frontend_covSum(Frontend_covSum), 	//Jaewon_regstate
	.Checking_Frontend_covmap(Frontend_covmap), 	//Jaewon_regstate
    .gated_clock(frontend_gated_clock),
    .reset(frontend_reset),
    .auto_icache_master_out_a_ready(frontend_auto_icache_master_out_a_ready),
    .auto_icache_master_out_a_valid(frontend_auto_icache_master_out_a_valid),
    .auto_icache_master_out_a_bits_address(frontend_auto_icache_master_out_a_bits_address),
    .auto_icache_master_out_d_valid(frontend_auto_icache_master_out_d_valid),
    .auto_icache_master_out_d_bits_opcode(frontend_auto_icache_master_out_d_bits_opcode),
    .auto_icache_master_out_d_bits_size(frontend_auto_icache_master_out_d_bits_size),
    .auto_icache_master_out_d_bits_data(frontend_auto_icache_master_out_d_bits_data),
    .auto_icache_master_out_d_bits_corrupt(frontend_auto_icache_master_out_d_bits_corrupt),
    .auto_reset_vector_sink_in(frontend_auto_reset_vector_sink_in),
    .io_cpu_might_request(frontend_io_cpu_might_request),
    .io_cpu_req_valid(frontend_io_cpu_req_valid),
    .io_cpu_req_bits_pc(frontend_io_cpu_req_bits_pc),
    .io_cpu_req_bits_speculative(frontend_io_cpu_req_bits_speculative),
    .io_cpu_sfence_valid(frontend_io_cpu_sfence_valid),
    .io_cpu_sfence_bits_rs1(frontend_io_cpu_sfence_bits_rs1),
    .io_cpu_sfence_bits_rs2(frontend_io_cpu_sfence_bits_rs2),
    .io_cpu_sfence_bits_addr(frontend_io_cpu_sfence_bits_addr),
    .io_cpu_resp_ready(frontend_io_cpu_resp_ready),
    .io_cpu_resp_valid(frontend_io_cpu_resp_valid),
    .io_cpu_resp_bits_btb_taken(frontend_io_cpu_resp_bits_btb_taken),
    .io_cpu_resp_bits_btb_bridx(frontend_io_cpu_resp_bits_btb_bridx),
    .io_cpu_resp_bits_btb_entry(frontend_io_cpu_resp_bits_btb_entry),
    .io_cpu_resp_bits_btb_bht_history(frontend_io_cpu_resp_bits_btb_bht_history),
    .io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_data(frontend_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_xcpt_pf_inst(frontend_io_cpu_resp_bits_xcpt_pf_inst),
    .io_cpu_resp_bits_xcpt_ae_inst(frontend_io_cpu_resp_bits_xcpt_ae_inst),
    .io_cpu_resp_bits_replay(frontend_io_cpu_resp_bits_replay),
    .io_cpu_btb_update_valid(frontend_io_cpu_btb_update_valid),
    .io_cpu_btb_update_bits_prediction_entry(frontend_io_cpu_btb_update_bits_prediction_entry),
    .io_cpu_btb_update_bits_pc(frontend_io_cpu_btb_update_bits_pc),
    .io_cpu_btb_update_bits_isValid(frontend_io_cpu_btb_update_bits_isValid),
    .io_cpu_btb_update_bits_br_pc(frontend_io_cpu_btb_update_bits_br_pc),
    .io_cpu_btb_update_bits_cfiType(frontend_io_cpu_btb_update_bits_cfiType),
    .io_cpu_bht_update_valid(frontend_io_cpu_bht_update_valid),
    .io_cpu_bht_update_bits_prediction_history(frontend_io_cpu_bht_update_bits_prediction_history),
    .io_cpu_bht_update_bits_pc(frontend_io_cpu_bht_update_bits_pc),
    .io_cpu_bht_update_bits_branch(frontend_io_cpu_bht_update_bits_branch),
    .io_cpu_bht_update_bits_taken(frontend_io_cpu_bht_update_bits_taken),
    .io_cpu_bht_update_bits_mispredict(frontend_io_cpu_bht_update_bits_mispredict),
    .io_cpu_flush_icache(frontend_io_cpu_flush_icache),
    .io_cpu_npc(frontend_io_cpu_npc),
    .io_ptw_req_ready(frontend_io_ptw_req_ready),
    .io_ptw_req_valid(frontend_io_ptw_req_valid),
    .io_ptw_req_bits_valid(frontend_io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr(frontend_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(frontend_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(frontend_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(frontend_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(frontend_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(frontend_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(frontend_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(frontend_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(frontend_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(frontend_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(frontend_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(frontend_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(frontend_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(frontend_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(frontend_io_ptw_ptbr_mode),
    .io_ptw_status_debug(frontend_io_ptw_status_debug),
    .io_ptw_status_prv(frontend_io_ptw_status_prv),
    .io_ptw_pmp_0_cfg_l(frontend_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(frontend_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(frontend_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(frontend_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(frontend_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(frontend_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(frontend_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(frontend_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(frontend_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(frontend_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(frontend_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(frontend_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(frontend_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(frontend_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(frontend_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(frontend_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(frontend_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(frontend_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(frontend_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(frontend_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(frontend_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(frontend_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(frontend_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(frontend_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(frontend_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(frontend_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(frontend_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(frontend_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(frontend_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(frontend_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(frontend_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(frontend_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(frontend_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(frontend_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(frontend_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(frontend_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(frontend_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(frontend_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(frontend_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(frontend_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(frontend_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(frontend_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(frontend_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(frontend_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(frontend_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(frontend_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(frontend_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(frontend_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(frontend_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(frontend_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(frontend_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(frontend_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(frontend_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(frontend_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(frontend_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(frontend_io_ptw_pmp_7_mask),
    .io_ptw_customCSRs_csrs_0_value(frontend_io_ptw_customCSRs_csrs_0_value),
    .io_covSum(frontend_io_covSum),
    .metaAssert(frontend_metaAssert),
    .metaReset(frontend_metaReset),
    .icache_halt(frontend_icache_halt),
    .fq_halt(frontend_fq_halt),
    .tlb_halt(frontend_tlb_halt),
    .btb_halt(frontend_btb_halt)
  );
  TLBuffer_7 buffer ( // @[Buffer.scala 69:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
    .auto_in_b_ready(buffer_auto_in_b_ready),
    .auto_in_b_valid(buffer_auto_in_b_valid),
    .auto_in_b_bits_opcode(buffer_auto_in_b_bits_opcode),
    .auto_in_b_bits_param(buffer_auto_in_b_bits_param),
    .auto_in_b_bits_size(buffer_auto_in_b_bits_size),
    .auto_in_b_bits_source(buffer_auto_in_b_bits_source),
    .auto_in_b_bits_address(buffer_auto_in_b_bits_address),
    .auto_in_b_bits_mask(buffer_auto_in_b_bits_mask),
    .auto_in_b_bits_corrupt(buffer_auto_in_b_bits_corrupt),
    .auto_in_c_ready(buffer_auto_in_c_ready),
    .auto_in_c_valid(buffer_auto_in_c_valid),
    .auto_in_c_bits_opcode(buffer_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(buffer_auto_in_c_bits_param),
    .auto_in_c_bits_size(buffer_auto_in_c_bits_size),
    .auto_in_c_bits_source(buffer_auto_in_c_bits_source),
    .auto_in_c_bits_address(buffer_auto_in_c_bits_address),
    .auto_in_c_bits_data(buffer_auto_in_c_bits_data),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_in_e_ready(buffer_auto_in_e_ready),
    .auto_in_e_valid(buffer_auto_in_e_valid),
    .auto_in_e_bits_sink(buffer_auto_in_e_bits_sink),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
    .auto_out_b_ready(buffer_auto_out_b_ready),
    .auto_out_b_valid(buffer_auto_out_b_valid),
    .auto_out_b_bits_opcode(buffer_auto_out_b_bits_opcode),
    .auto_out_b_bits_param(buffer_auto_out_b_bits_param),
    .auto_out_b_bits_size(buffer_auto_out_b_bits_size),
    .auto_out_b_bits_source(buffer_auto_out_b_bits_source),
    .auto_out_b_bits_address(buffer_auto_out_b_bits_address),
    .auto_out_b_bits_mask(buffer_auto_out_b_bits_mask),
    .auto_out_b_bits_corrupt(buffer_auto_out_b_bits_corrupt),
    .auto_out_c_ready(buffer_auto_out_c_ready),
    .auto_out_c_valid(buffer_auto_out_c_valid),
    .auto_out_c_bits_opcode(buffer_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(buffer_auto_out_c_bits_param),
    .auto_out_c_bits_size(buffer_auto_out_c_bits_size),
    .auto_out_c_bits_source(buffer_auto_out_c_bits_source),
    .auto_out_c_bits_address(buffer_auto_out_c_bits_address),
    .auto_out_c_bits_data(buffer_auto_out_c_bits_data),
    .auto_out_c_bits_corrupt(buffer_auto_out_c_bits_corrupt),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(buffer_auto_out_d_bits_param),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_sink(buffer_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt),
    .auto_out_e_ready(buffer_auto_out_e_ready),
    .auto_out_e_valid(buffer_auto_out_e_valid),
    .auto_out_e_bits_sink(buffer_auto_out_e_bits_sink),
    .io_covSum(buffer_io_covSum),
    .metaAssert(buffer_metaAssert),
    .metaReset(buffer_metaReset),
    .Queue_3_halt(buffer_Queue_3_halt),
    .Queue_halt(buffer_Queue_halt),
    .TLMonitor_halt(buffer_TLMonitor_halt),
    .Queue_2_halt(buffer_Queue_2_halt),
    .Queue_4_halt(buffer_Queue_4_halt),
    .Queue_1_halt(buffer_Queue_1_halt)
  );
  IntSyncAsyncCrossingSink intsink ( // @[Crossing.scala 74:29]
    .clock(intsink_clock),
    .auto_in_sync_0(intsink_auto_in_sync_0),
    .auto_out_0(intsink_auto_out_0),
    .io_covSum(intsink_io_covSum),
    .metaAssert(intsink_metaAssert),
    .metaReset(intsink_metaReset),
    .SynchronizerShiftReg_w1_d3_halt(intsink_SynchronizerShiftReg_w1_d3_halt)
  );
  IntSyncSyncCrossingSink intsink_1 ( // @[Crossing.scala 94:29]
    .auto_in_sync_0(intsink_1_auto_in_sync_0),
    .auto_in_sync_1(intsink_1_auto_in_sync_1),
    .auto_out_0(intsink_1_auto_out_0),
    .auto_out_1(intsink_1_auto_out_1),
    .io_covSum(intsink_1_io_covSum),
    .metaAssert(intsink_1_metaAssert)
  );
  IntSyncSyncCrossingSink_1 intsink_2 ( // @[Crossing.scala 94:29]
    .auto_in_sync_0(intsink_2_auto_in_sync_0),
    .auto_out_0(intsink_2_auto_out_0),
    .io_covSum(intsink_2_io_covSum),
    .metaAssert(intsink_2_metaAssert)
  );
  IntSyncSyncCrossingSink_1 intsink_3 ( // @[Crossing.scala 94:29]
    .auto_in_sync_0(intsink_3_auto_in_sync_0),
    .auto_out_0(intsink_3_auto_out_0),
    .io_covSum(intsink_3_io_covSum),
    .metaAssert(intsink_3_metaAssert)
  );
  FPU fpuOpt ( // @[RocketTile.scala 195:62]
    .clock(fpuOpt_clock),
    .reset(fpuOpt_reset),
    .io_inst(fpuOpt_io_inst),
    .io_fromint_data(fpuOpt_io_fromint_data),
    .io_fcsr_rm(fpuOpt_io_fcsr_rm),
    .io_fcsr_flags_valid(fpuOpt_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(fpuOpt_io_fcsr_flags_bits),
    .io_store_data(fpuOpt_io_store_data),
    .io_toint_data(fpuOpt_io_toint_data),
    .io_dmem_resp_val(fpuOpt_io_dmem_resp_val),
    .io_dmem_resp_type(fpuOpt_io_dmem_resp_type),
    .io_dmem_resp_tag(fpuOpt_io_dmem_resp_tag),
    .io_dmem_resp_data(fpuOpt_io_dmem_resp_data),
    .io_valid(fpuOpt_io_valid),
    .io_fcsr_rdy(fpuOpt_io_fcsr_rdy),
    .io_nack_mem(fpuOpt_io_nack_mem),
    .io_illegal_rm(fpuOpt_io_illegal_rm),
    .io_killx(fpuOpt_io_killx),
    .io_killm(fpuOpt_io_killm),
    .io_dec_wen(fpuOpt_io_dec_wen),
    .io_dec_ren1(fpuOpt_io_dec_ren1),
    .io_dec_ren2(fpuOpt_io_dec_ren2),
    .io_dec_ren3(fpuOpt_io_dec_ren3),
    .io_sboard_set(fpuOpt_io_sboard_set),
    .io_sboard_clr(fpuOpt_io_sboard_clr),
    .io_sboard_clra(fpuOpt_io_sboard_clra),
    .io_covSum(fpuOpt_io_covSum),
    .metaAssert(fpuOpt_metaAssert),
    .metaReset(fpuOpt_metaReset),
    .divSqrt_1_halt(fpuOpt_divSqrt_1_halt),
    .ifpu_halt(fpuOpt_ifpu_halt),
    .divSqrt_halt(fpuOpt_divSqrt_halt),
    .fpmu_halt(fpuOpt_fpmu_halt),
    .dfma_halt(fpuOpt_dfma_halt),
    .fpiu_halt(fpuOpt_fpiu_halt),
    .sfma_halt(fpuOpt_sfma_halt),
    .Checking_FPU_regstate(FPU_regstate),		//Jaewon_FPU_regstate
    .Checking_FPU_covSum(FPU_covSum)		   //Jaewon_FPU_regstate
  );
  HellaCacheArbiter dcacheArb ( // @[HellaCache.scala 264:25]
    .clock(dcacheArb_clock),
    .io_requestor_0_req_ready(dcacheArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dcacheArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(dcacheArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_s1_kill(dcacheArb_io_requestor_0_s1_kill),
    .io_requestor_0_s2_nack(dcacheArb_io_requestor_0_s2_nack),
    .io_requestor_0_resp_valid(dcacheArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_data(dcacheArb_io_requestor_0_resp_bits_data),
    .io_requestor_0_s2_xcpt_ae_ld(dcacheArb_io_requestor_0_s2_xcpt_ae_ld),
    .io_requestor_1_req_ready(dcacheArb_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(dcacheArb_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(dcacheArb_io_requestor_1_req_bits_addr),
    .io_requestor_1_req_bits_tag(dcacheArb_io_requestor_1_req_bits_tag),
    .io_requestor_1_req_bits_cmd(dcacheArb_io_requestor_1_req_bits_cmd),
    .io_requestor_1_req_bits_size(dcacheArb_io_requestor_1_req_bits_size),
    .io_requestor_1_req_bits_signed(dcacheArb_io_requestor_1_req_bits_signed),
    .io_requestor_1_s1_kill(dcacheArb_io_requestor_1_s1_kill),
    .io_requestor_1_s1_data_data(dcacheArb_io_requestor_1_s1_data_data),
    .io_requestor_1_s2_nack(dcacheArb_io_requestor_1_s2_nack),
    .io_requestor_1_resp_valid(dcacheArb_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_tag(dcacheArb_io_requestor_1_resp_bits_tag),
    .io_requestor_1_resp_bits_size(dcacheArb_io_requestor_1_resp_bits_size),
    .io_requestor_1_resp_bits_data(dcacheArb_io_requestor_1_resp_bits_data),
    .io_requestor_1_resp_bits_replay(dcacheArb_io_requestor_1_resp_bits_replay),
    .io_requestor_1_resp_bits_has_data(dcacheArb_io_requestor_1_resp_bits_has_data),
    .io_requestor_1_resp_bits_data_word_bypass(dcacheArb_io_requestor_1_resp_bits_data_word_bypass),
    .io_requestor_1_replay_next(dcacheArb_io_requestor_1_replay_next),
    .io_requestor_1_s2_xcpt_ma_ld(dcacheArb_io_requestor_1_s2_xcpt_ma_ld),
    .io_requestor_1_s2_xcpt_ma_st(dcacheArb_io_requestor_1_s2_xcpt_ma_st),
    .io_requestor_1_s2_xcpt_pf_ld(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),
    .io_requestor_1_s2_xcpt_pf_st(dcacheArb_io_requestor_1_s2_xcpt_pf_st),
    .io_requestor_1_s2_xcpt_ae_ld(dcacheArb_io_requestor_1_s2_xcpt_ae_ld),
    .io_requestor_1_s2_xcpt_ae_st(dcacheArb_io_requestor_1_s2_xcpt_ae_st),
    .io_requestor_1_ordered(dcacheArb_io_requestor_1_ordered),
    .io_requestor_1_perf_release(dcacheArb_io_requestor_1_perf_release),
    .io_requestor_1_perf_grant(dcacheArb_io_requestor_1_perf_grant),
    .io_mem_req_ready(dcacheArb_io_mem_req_ready),
    .io_mem_req_valid(dcacheArb_io_mem_req_valid),
    .io_mem_req_bits_addr(dcacheArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(dcacheArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(dcacheArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_size(dcacheArb_io_mem_req_bits_size),
    .io_mem_req_bits_signed(dcacheArb_io_mem_req_bits_signed),
    .io_mem_req_bits_phys(dcacheArb_io_mem_req_bits_phys),
    .io_mem_s1_kill(dcacheArb_io_mem_s1_kill),
    .io_mem_s1_data_data(dcacheArb_io_mem_s1_data_data),
    .io_mem_s2_nack(dcacheArb_io_mem_s2_nack),
    .io_mem_resp_valid(dcacheArb_io_mem_resp_valid),
    .io_mem_resp_bits_tag(dcacheArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_size(dcacheArb_io_mem_resp_bits_size),
    .io_mem_resp_bits_data(dcacheArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(dcacheArb_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(dcacheArb_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(dcacheArb_io_mem_resp_bits_data_word_bypass),
    .io_mem_replay_next(dcacheArb_io_mem_replay_next),
    .io_mem_s2_xcpt_ma_ld(dcacheArb_io_mem_s2_xcpt_ma_ld),
    .io_mem_s2_xcpt_ma_st(dcacheArb_io_mem_s2_xcpt_ma_st),
    .io_mem_s2_xcpt_pf_ld(dcacheArb_io_mem_s2_xcpt_pf_ld),
    .io_mem_s2_xcpt_pf_st(dcacheArb_io_mem_s2_xcpt_pf_st),
    .io_mem_s2_xcpt_ae_ld(dcacheArb_io_mem_s2_xcpt_ae_ld),
    .io_mem_s2_xcpt_ae_st(dcacheArb_io_mem_s2_xcpt_ae_st),
    .io_mem_ordered(dcacheArb_io_mem_ordered),
    .io_mem_perf_release(dcacheArb_io_mem_perf_release),
    .io_mem_perf_grant(dcacheArb_io_mem_perf_grant),
    .io_covSum(dcacheArb_io_covSum),
    .metaAssert(dcacheArb_metaAssert),
    .metaReset(dcacheArb_metaReset)
  );
  PTW ptw ( // @[PTW.scala 395:19]
    .clock(ptw_clock),
    .reset(ptw_reset),
    .io_requestor_0_req_ready(ptw_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(ptw_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_bits_addr(ptw_io_requestor_0_req_bits_bits_addr),
    .io_requestor_0_resp_valid(ptw_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_ae(ptw_io_requestor_0_resp_bits_ae),
    .io_requestor_0_resp_bits_pte_ppn(ptw_io_requestor_0_resp_bits_pte_ppn),
    .io_requestor_0_resp_bits_pte_d(ptw_io_requestor_0_resp_bits_pte_d),
    .io_requestor_0_resp_bits_pte_a(ptw_io_requestor_0_resp_bits_pte_a),
    .io_requestor_0_resp_bits_pte_g(ptw_io_requestor_0_resp_bits_pte_g),
    .io_requestor_0_resp_bits_pte_u(ptw_io_requestor_0_resp_bits_pte_u),
    .io_requestor_0_resp_bits_pte_x(ptw_io_requestor_0_resp_bits_pte_x),
    .io_requestor_0_resp_bits_pte_w(ptw_io_requestor_0_resp_bits_pte_w),
    .io_requestor_0_resp_bits_pte_r(ptw_io_requestor_0_resp_bits_pte_r),
    .io_requestor_0_resp_bits_pte_v(ptw_io_requestor_0_resp_bits_pte_v),
    .io_requestor_0_resp_bits_level(ptw_io_requestor_0_resp_bits_level),
    .io_requestor_0_resp_bits_homogeneous(ptw_io_requestor_0_resp_bits_homogeneous),
    .io_requestor_0_ptbr_mode(ptw_io_requestor_0_ptbr_mode),
    .io_requestor_0_status_debug(ptw_io_requestor_0_status_debug),
    .io_requestor_0_status_dprv(ptw_io_requestor_0_status_dprv),
    .io_requestor_0_status_mxr(ptw_io_requestor_0_status_mxr),
    .io_requestor_0_status_sum(ptw_io_requestor_0_status_sum),
    .io_requestor_0_pmp_0_cfg_l(ptw_io_requestor_0_pmp_0_cfg_l),
    .io_requestor_0_pmp_0_cfg_a(ptw_io_requestor_0_pmp_0_cfg_a),
    .io_requestor_0_pmp_0_cfg_x(ptw_io_requestor_0_pmp_0_cfg_x),
    .io_requestor_0_pmp_0_cfg_w(ptw_io_requestor_0_pmp_0_cfg_w),
    .io_requestor_0_pmp_0_cfg_r(ptw_io_requestor_0_pmp_0_cfg_r),
    .io_requestor_0_pmp_0_addr(ptw_io_requestor_0_pmp_0_addr),
    .io_requestor_0_pmp_0_mask(ptw_io_requestor_0_pmp_0_mask),
    .io_requestor_0_pmp_1_cfg_l(ptw_io_requestor_0_pmp_1_cfg_l),
    .io_requestor_0_pmp_1_cfg_a(ptw_io_requestor_0_pmp_1_cfg_a),
    .io_requestor_0_pmp_1_cfg_x(ptw_io_requestor_0_pmp_1_cfg_x),
    .io_requestor_0_pmp_1_cfg_w(ptw_io_requestor_0_pmp_1_cfg_w),
    .io_requestor_0_pmp_1_cfg_r(ptw_io_requestor_0_pmp_1_cfg_r),
    .io_requestor_0_pmp_1_addr(ptw_io_requestor_0_pmp_1_addr),
    .io_requestor_0_pmp_1_mask(ptw_io_requestor_0_pmp_1_mask),
    .io_requestor_0_pmp_2_cfg_l(ptw_io_requestor_0_pmp_2_cfg_l),
    .io_requestor_0_pmp_2_cfg_a(ptw_io_requestor_0_pmp_2_cfg_a),
    .io_requestor_0_pmp_2_cfg_x(ptw_io_requestor_0_pmp_2_cfg_x),
    .io_requestor_0_pmp_2_cfg_w(ptw_io_requestor_0_pmp_2_cfg_w),
    .io_requestor_0_pmp_2_cfg_r(ptw_io_requestor_0_pmp_2_cfg_r),
    .io_requestor_0_pmp_2_addr(ptw_io_requestor_0_pmp_2_addr),
    .io_requestor_0_pmp_2_mask(ptw_io_requestor_0_pmp_2_mask),
    .io_requestor_0_pmp_3_cfg_l(ptw_io_requestor_0_pmp_3_cfg_l),
    .io_requestor_0_pmp_3_cfg_a(ptw_io_requestor_0_pmp_3_cfg_a),
    .io_requestor_0_pmp_3_cfg_x(ptw_io_requestor_0_pmp_3_cfg_x),
    .io_requestor_0_pmp_3_cfg_w(ptw_io_requestor_0_pmp_3_cfg_w),
    .io_requestor_0_pmp_3_cfg_r(ptw_io_requestor_0_pmp_3_cfg_r),
    .io_requestor_0_pmp_3_addr(ptw_io_requestor_0_pmp_3_addr),
    .io_requestor_0_pmp_3_mask(ptw_io_requestor_0_pmp_3_mask),
    .io_requestor_0_pmp_4_cfg_l(ptw_io_requestor_0_pmp_4_cfg_l),
    .io_requestor_0_pmp_4_cfg_a(ptw_io_requestor_0_pmp_4_cfg_a),
    .io_requestor_0_pmp_4_cfg_x(ptw_io_requestor_0_pmp_4_cfg_x),
    .io_requestor_0_pmp_4_cfg_w(ptw_io_requestor_0_pmp_4_cfg_w),
    .io_requestor_0_pmp_4_cfg_r(ptw_io_requestor_0_pmp_4_cfg_r),
    .io_requestor_0_pmp_4_addr(ptw_io_requestor_0_pmp_4_addr),
    .io_requestor_0_pmp_4_mask(ptw_io_requestor_0_pmp_4_mask),
    .io_requestor_0_pmp_5_cfg_l(ptw_io_requestor_0_pmp_5_cfg_l),
    .io_requestor_0_pmp_5_cfg_a(ptw_io_requestor_0_pmp_5_cfg_a),
    .io_requestor_0_pmp_5_cfg_x(ptw_io_requestor_0_pmp_5_cfg_x),
    .io_requestor_0_pmp_5_cfg_w(ptw_io_requestor_0_pmp_5_cfg_w),
    .io_requestor_0_pmp_5_cfg_r(ptw_io_requestor_0_pmp_5_cfg_r),
    .io_requestor_0_pmp_5_addr(ptw_io_requestor_0_pmp_5_addr),
    .io_requestor_0_pmp_5_mask(ptw_io_requestor_0_pmp_5_mask),
    .io_requestor_0_pmp_6_cfg_l(ptw_io_requestor_0_pmp_6_cfg_l),
    .io_requestor_0_pmp_6_cfg_a(ptw_io_requestor_0_pmp_6_cfg_a),
    .io_requestor_0_pmp_6_cfg_x(ptw_io_requestor_0_pmp_6_cfg_x),
    .io_requestor_0_pmp_6_cfg_w(ptw_io_requestor_0_pmp_6_cfg_w),
    .io_requestor_0_pmp_6_cfg_r(ptw_io_requestor_0_pmp_6_cfg_r),
    .io_requestor_0_pmp_6_addr(ptw_io_requestor_0_pmp_6_addr),
    .io_requestor_0_pmp_6_mask(ptw_io_requestor_0_pmp_6_mask),
    .io_requestor_0_pmp_7_cfg_l(ptw_io_requestor_0_pmp_7_cfg_l),
    .io_requestor_0_pmp_7_cfg_a(ptw_io_requestor_0_pmp_7_cfg_a),
    .io_requestor_0_pmp_7_cfg_x(ptw_io_requestor_0_pmp_7_cfg_x),
    .io_requestor_0_pmp_7_cfg_w(ptw_io_requestor_0_pmp_7_cfg_w),
    .io_requestor_0_pmp_7_cfg_r(ptw_io_requestor_0_pmp_7_cfg_r),
    .io_requestor_0_pmp_7_addr(ptw_io_requestor_0_pmp_7_addr),
    .io_requestor_0_pmp_7_mask(ptw_io_requestor_0_pmp_7_mask),
    .io_requestor_1_req_ready(ptw_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(ptw_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_valid(ptw_io_requestor_1_req_bits_valid),
    .io_requestor_1_req_bits_bits_addr(ptw_io_requestor_1_req_bits_bits_addr),
    .io_requestor_1_resp_valid(ptw_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_ae(ptw_io_requestor_1_resp_bits_ae),
    .io_requestor_1_resp_bits_pte_ppn(ptw_io_requestor_1_resp_bits_pte_ppn),
    .io_requestor_1_resp_bits_pte_d(ptw_io_requestor_1_resp_bits_pte_d),
    .io_requestor_1_resp_bits_pte_a(ptw_io_requestor_1_resp_bits_pte_a),
    .io_requestor_1_resp_bits_pte_g(ptw_io_requestor_1_resp_bits_pte_g),
    .io_requestor_1_resp_bits_pte_u(ptw_io_requestor_1_resp_bits_pte_u),
    .io_requestor_1_resp_bits_pte_x(ptw_io_requestor_1_resp_bits_pte_x),
    .io_requestor_1_resp_bits_pte_w(ptw_io_requestor_1_resp_bits_pte_w),
    .io_requestor_1_resp_bits_pte_r(ptw_io_requestor_1_resp_bits_pte_r),
    .io_requestor_1_resp_bits_pte_v(ptw_io_requestor_1_resp_bits_pte_v),
    .io_requestor_1_resp_bits_level(ptw_io_requestor_1_resp_bits_level),
    .io_requestor_1_resp_bits_homogeneous(ptw_io_requestor_1_resp_bits_homogeneous),
    .io_requestor_1_ptbr_mode(ptw_io_requestor_1_ptbr_mode),
    .io_requestor_1_status_debug(ptw_io_requestor_1_status_debug),
    .io_requestor_1_status_prv(ptw_io_requestor_1_status_prv),
    .io_requestor_1_pmp_0_cfg_l(ptw_io_requestor_1_pmp_0_cfg_l),
    .io_requestor_1_pmp_0_cfg_a(ptw_io_requestor_1_pmp_0_cfg_a),
    .io_requestor_1_pmp_0_cfg_x(ptw_io_requestor_1_pmp_0_cfg_x),
    .io_requestor_1_pmp_0_cfg_w(ptw_io_requestor_1_pmp_0_cfg_w),
    .io_requestor_1_pmp_0_cfg_r(ptw_io_requestor_1_pmp_0_cfg_r),
    .io_requestor_1_pmp_0_addr(ptw_io_requestor_1_pmp_0_addr),
    .io_requestor_1_pmp_0_mask(ptw_io_requestor_1_pmp_0_mask),
    .io_requestor_1_pmp_1_cfg_l(ptw_io_requestor_1_pmp_1_cfg_l),
    .io_requestor_1_pmp_1_cfg_a(ptw_io_requestor_1_pmp_1_cfg_a),
    .io_requestor_1_pmp_1_cfg_x(ptw_io_requestor_1_pmp_1_cfg_x),
    .io_requestor_1_pmp_1_cfg_w(ptw_io_requestor_1_pmp_1_cfg_w),
    .io_requestor_1_pmp_1_cfg_r(ptw_io_requestor_1_pmp_1_cfg_r),
    .io_requestor_1_pmp_1_addr(ptw_io_requestor_1_pmp_1_addr),
    .io_requestor_1_pmp_1_mask(ptw_io_requestor_1_pmp_1_mask),
    .io_requestor_1_pmp_2_cfg_l(ptw_io_requestor_1_pmp_2_cfg_l),
    .io_requestor_1_pmp_2_cfg_a(ptw_io_requestor_1_pmp_2_cfg_a),
    .io_requestor_1_pmp_2_cfg_x(ptw_io_requestor_1_pmp_2_cfg_x),
    .io_requestor_1_pmp_2_cfg_w(ptw_io_requestor_1_pmp_2_cfg_w),
    .io_requestor_1_pmp_2_cfg_r(ptw_io_requestor_1_pmp_2_cfg_r),
    .io_requestor_1_pmp_2_addr(ptw_io_requestor_1_pmp_2_addr),
    .io_requestor_1_pmp_2_mask(ptw_io_requestor_1_pmp_2_mask),
    .io_requestor_1_pmp_3_cfg_l(ptw_io_requestor_1_pmp_3_cfg_l),
    .io_requestor_1_pmp_3_cfg_a(ptw_io_requestor_1_pmp_3_cfg_a),
    .io_requestor_1_pmp_3_cfg_x(ptw_io_requestor_1_pmp_3_cfg_x),
    .io_requestor_1_pmp_3_cfg_w(ptw_io_requestor_1_pmp_3_cfg_w),
    .io_requestor_1_pmp_3_cfg_r(ptw_io_requestor_1_pmp_3_cfg_r),
    .io_requestor_1_pmp_3_addr(ptw_io_requestor_1_pmp_3_addr),
    .io_requestor_1_pmp_3_mask(ptw_io_requestor_1_pmp_3_mask),
    .io_requestor_1_pmp_4_cfg_l(ptw_io_requestor_1_pmp_4_cfg_l),
    .io_requestor_1_pmp_4_cfg_a(ptw_io_requestor_1_pmp_4_cfg_a),
    .io_requestor_1_pmp_4_cfg_x(ptw_io_requestor_1_pmp_4_cfg_x),
    .io_requestor_1_pmp_4_cfg_w(ptw_io_requestor_1_pmp_4_cfg_w),
    .io_requestor_1_pmp_4_cfg_r(ptw_io_requestor_1_pmp_4_cfg_r),
    .io_requestor_1_pmp_4_addr(ptw_io_requestor_1_pmp_4_addr),
    .io_requestor_1_pmp_4_mask(ptw_io_requestor_1_pmp_4_mask),
    .io_requestor_1_pmp_5_cfg_l(ptw_io_requestor_1_pmp_5_cfg_l),
    .io_requestor_1_pmp_5_cfg_a(ptw_io_requestor_1_pmp_5_cfg_a),
    .io_requestor_1_pmp_5_cfg_x(ptw_io_requestor_1_pmp_5_cfg_x),
    .io_requestor_1_pmp_5_cfg_w(ptw_io_requestor_1_pmp_5_cfg_w),
    .io_requestor_1_pmp_5_cfg_r(ptw_io_requestor_1_pmp_5_cfg_r),
    .io_requestor_1_pmp_5_addr(ptw_io_requestor_1_pmp_5_addr),
    .io_requestor_1_pmp_5_mask(ptw_io_requestor_1_pmp_5_mask),
    .io_requestor_1_pmp_6_cfg_l(ptw_io_requestor_1_pmp_6_cfg_l),
    .io_requestor_1_pmp_6_cfg_a(ptw_io_requestor_1_pmp_6_cfg_a),
    .io_requestor_1_pmp_6_cfg_x(ptw_io_requestor_1_pmp_6_cfg_x),
    .io_requestor_1_pmp_6_cfg_w(ptw_io_requestor_1_pmp_6_cfg_w),
    .io_requestor_1_pmp_6_cfg_r(ptw_io_requestor_1_pmp_6_cfg_r),
    .io_requestor_1_pmp_6_addr(ptw_io_requestor_1_pmp_6_addr),
    .io_requestor_1_pmp_6_mask(ptw_io_requestor_1_pmp_6_mask),
    .io_requestor_1_pmp_7_cfg_l(ptw_io_requestor_1_pmp_7_cfg_l),
    .io_requestor_1_pmp_7_cfg_a(ptw_io_requestor_1_pmp_7_cfg_a),
    .io_requestor_1_pmp_7_cfg_x(ptw_io_requestor_1_pmp_7_cfg_x),
    .io_requestor_1_pmp_7_cfg_w(ptw_io_requestor_1_pmp_7_cfg_w),
    .io_requestor_1_pmp_7_cfg_r(ptw_io_requestor_1_pmp_7_cfg_r),
    .io_requestor_1_pmp_7_addr(ptw_io_requestor_1_pmp_7_addr),
    .io_requestor_1_pmp_7_mask(ptw_io_requestor_1_pmp_7_mask),
    .io_requestor_1_customCSRs_csrs_0_value(ptw_io_requestor_1_customCSRs_csrs_0_value),
    .io_mem_req_ready(ptw_io_mem_req_ready),
    .io_mem_req_valid(ptw_io_mem_req_valid),
    .io_mem_req_bits_addr(ptw_io_mem_req_bits_addr),
    .io_mem_s1_kill(ptw_io_mem_s1_kill),
    .io_mem_s2_nack(ptw_io_mem_s2_nack),
    .io_mem_resp_valid(ptw_io_mem_resp_valid),
    .io_mem_resp_bits_data(ptw_io_mem_resp_bits_data),
    .io_mem_s2_xcpt_ae_ld(ptw_io_mem_s2_xcpt_ae_ld),
    .io_dpath_ptbr_mode(ptw_io_dpath_ptbr_mode),
    .io_dpath_ptbr_ppn(ptw_io_dpath_ptbr_ppn),
    .io_dpath_sfence_valid(ptw_io_dpath_sfence_valid),
    .io_dpath_sfence_bits_rs1(ptw_io_dpath_sfence_bits_rs1),
    .io_dpath_status_debug(ptw_io_dpath_status_debug),
    .io_dpath_status_dprv(ptw_io_dpath_status_dprv),
    .io_dpath_status_prv(ptw_io_dpath_status_prv),
    .io_dpath_status_mxr(ptw_io_dpath_status_mxr),
    .io_dpath_status_sum(ptw_io_dpath_status_sum),
    .io_dpath_pmp_0_cfg_l(ptw_io_dpath_pmp_0_cfg_l),
    .io_dpath_pmp_0_cfg_a(ptw_io_dpath_pmp_0_cfg_a),
    .io_dpath_pmp_0_cfg_x(ptw_io_dpath_pmp_0_cfg_x),
    .io_dpath_pmp_0_cfg_w(ptw_io_dpath_pmp_0_cfg_w),
    .io_dpath_pmp_0_cfg_r(ptw_io_dpath_pmp_0_cfg_r),
    .io_dpath_pmp_0_addr(ptw_io_dpath_pmp_0_addr),
    .io_dpath_pmp_0_mask(ptw_io_dpath_pmp_0_mask),
    .io_dpath_pmp_1_cfg_l(ptw_io_dpath_pmp_1_cfg_l),
    .io_dpath_pmp_1_cfg_a(ptw_io_dpath_pmp_1_cfg_a),
    .io_dpath_pmp_1_cfg_x(ptw_io_dpath_pmp_1_cfg_x),
    .io_dpath_pmp_1_cfg_w(ptw_io_dpath_pmp_1_cfg_w),
    .io_dpath_pmp_1_cfg_r(ptw_io_dpath_pmp_1_cfg_r),
    .io_dpath_pmp_1_addr(ptw_io_dpath_pmp_1_addr),
    .io_dpath_pmp_1_mask(ptw_io_dpath_pmp_1_mask),
    .io_dpath_pmp_2_cfg_l(ptw_io_dpath_pmp_2_cfg_l),
    .io_dpath_pmp_2_cfg_a(ptw_io_dpath_pmp_2_cfg_a),
    .io_dpath_pmp_2_cfg_x(ptw_io_dpath_pmp_2_cfg_x),
    .io_dpath_pmp_2_cfg_w(ptw_io_dpath_pmp_2_cfg_w),
    .io_dpath_pmp_2_cfg_r(ptw_io_dpath_pmp_2_cfg_r),
    .io_dpath_pmp_2_addr(ptw_io_dpath_pmp_2_addr),
    .io_dpath_pmp_2_mask(ptw_io_dpath_pmp_2_mask),
    .io_dpath_pmp_3_cfg_l(ptw_io_dpath_pmp_3_cfg_l),
    .io_dpath_pmp_3_cfg_a(ptw_io_dpath_pmp_3_cfg_a),
    .io_dpath_pmp_3_cfg_x(ptw_io_dpath_pmp_3_cfg_x),
    .io_dpath_pmp_3_cfg_w(ptw_io_dpath_pmp_3_cfg_w),
    .io_dpath_pmp_3_cfg_r(ptw_io_dpath_pmp_3_cfg_r),
    .io_dpath_pmp_3_addr(ptw_io_dpath_pmp_3_addr),
    .io_dpath_pmp_3_mask(ptw_io_dpath_pmp_3_mask),
    .io_dpath_pmp_4_cfg_l(ptw_io_dpath_pmp_4_cfg_l),
    .io_dpath_pmp_4_cfg_a(ptw_io_dpath_pmp_4_cfg_a),
    .io_dpath_pmp_4_cfg_x(ptw_io_dpath_pmp_4_cfg_x),
    .io_dpath_pmp_4_cfg_w(ptw_io_dpath_pmp_4_cfg_w),
    .io_dpath_pmp_4_cfg_r(ptw_io_dpath_pmp_4_cfg_r),
    .io_dpath_pmp_4_addr(ptw_io_dpath_pmp_4_addr),
    .io_dpath_pmp_4_mask(ptw_io_dpath_pmp_4_mask),
    .io_dpath_pmp_5_cfg_l(ptw_io_dpath_pmp_5_cfg_l),
    .io_dpath_pmp_5_cfg_a(ptw_io_dpath_pmp_5_cfg_a),
    .io_dpath_pmp_5_cfg_x(ptw_io_dpath_pmp_5_cfg_x),
    .io_dpath_pmp_5_cfg_w(ptw_io_dpath_pmp_5_cfg_w),
    .io_dpath_pmp_5_cfg_r(ptw_io_dpath_pmp_5_cfg_r),
    .io_dpath_pmp_5_addr(ptw_io_dpath_pmp_5_addr),
    .io_dpath_pmp_5_mask(ptw_io_dpath_pmp_5_mask),
    .io_dpath_pmp_6_cfg_l(ptw_io_dpath_pmp_6_cfg_l),
    .io_dpath_pmp_6_cfg_a(ptw_io_dpath_pmp_6_cfg_a),
    .io_dpath_pmp_6_cfg_x(ptw_io_dpath_pmp_6_cfg_x),
    .io_dpath_pmp_6_cfg_w(ptw_io_dpath_pmp_6_cfg_w),
    .io_dpath_pmp_6_cfg_r(ptw_io_dpath_pmp_6_cfg_r),
    .io_dpath_pmp_6_addr(ptw_io_dpath_pmp_6_addr),
    .io_dpath_pmp_6_mask(ptw_io_dpath_pmp_6_mask),
    .io_dpath_pmp_7_cfg_l(ptw_io_dpath_pmp_7_cfg_l),
    .io_dpath_pmp_7_cfg_a(ptw_io_dpath_pmp_7_cfg_a),
    .io_dpath_pmp_7_cfg_x(ptw_io_dpath_pmp_7_cfg_x),
    .io_dpath_pmp_7_cfg_w(ptw_io_dpath_pmp_7_cfg_w),
    .io_dpath_pmp_7_cfg_r(ptw_io_dpath_pmp_7_cfg_r),
    .io_dpath_pmp_7_addr(ptw_io_dpath_pmp_7_addr),
    .io_dpath_pmp_7_mask(ptw_io_dpath_pmp_7_mask),
    .io_dpath_customCSRs_csrs_0_value(ptw_io_dpath_customCSRs_csrs_0_value),
    .io_covSum(ptw_io_covSum),
    .metaAssert(ptw_metaAssert),
    .metaReset(ptw_metaReset),
    .Checking_PTW_covSum(PTW_covSum),				//Jaewon_PTW_covSum
    .Checking_PTW_regstate(PTW_regstate)			//Jaewon_PTW_regstate
  );
  Rocket core ( // @[RocketTile.scala 135:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_hartid(core_io_hartid),
    .io_interrupts_debug(core_io_interrupts_debug),
    .io_interrupts_mtip(core_io_interrupts_mtip),
    .io_interrupts_msip(core_io_interrupts_msip),
    .io_interrupts_meip(core_io_interrupts_meip),
    .io_interrupts_seip(core_io_interrupts_seip),
    .io_imem_might_request(core_io_imem_might_request),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_pc(core_io_imem_req_bits_pc),
    .io_imem_req_bits_speculative(core_io_imem_req_bits_speculative),
    .io_imem_sfence_valid(core_io_imem_sfence_valid),
    .io_imem_sfence_bits_rs1(core_io_imem_sfence_bits_rs1),
    .io_imem_sfence_bits_rs2(core_io_imem_sfence_bits_rs2),
    .io_imem_sfence_bits_addr(core_io_imem_sfence_bits_addr),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_btb_taken(core_io_imem_resp_bits_btb_taken),
    .io_imem_resp_bits_btb_bridx(core_io_imem_resp_bits_btb_bridx),
    .io_imem_resp_bits_btb_entry(core_io_imem_resp_bits_btb_entry),
    .io_imem_resp_bits_btb_bht_history(core_io_imem_resp_bits_btb_bht_history),
    .io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data(core_io_imem_resp_bits_data),
    .io_imem_resp_bits_xcpt_pf_inst(core_io_imem_resp_bits_xcpt_pf_inst),
    .io_imem_resp_bits_xcpt_ae_inst(core_io_imem_resp_bits_xcpt_ae_inst),
    .io_imem_resp_bits_replay(core_io_imem_resp_bits_replay),
    .io_imem_btb_update_valid(core_io_imem_btb_update_valid),
    .io_imem_btb_update_bits_prediction_entry(core_io_imem_btb_update_bits_prediction_entry),
    .io_imem_btb_update_bits_pc(core_io_imem_btb_update_bits_pc),
    .io_imem_btb_update_bits_isValid(core_io_imem_btb_update_bits_isValid),
    .io_imem_btb_update_bits_br_pc(core_io_imem_btb_update_bits_br_pc),
    .io_imem_btb_update_bits_cfiType(core_io_imem_btb_update_bits_cfiType),
    .io_imem_bht_update_valid(core_io_imem_bht_update_valid),
    .io_imem_bht_update_bits_prediction_history(core_io_imem_bht_update_bits_prediction_history),
    .io_imem_bht_update_bits_pc(core_io_imem_bht_update_bits_pc),
    .io_imem_bht_update_bits_branch(core_io_imem_bht_update_bits_branch),
    .io_imem_bht_update_bits_taken(core_io_imem_bht_update_bits_taken),
    .io_imem_bht_update_bits_mispredict(core_io_imem_bht_update_bits_mispredict),
    .io_imem_flush_icache(core_io_imem_flush_icache),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_size(core_io_dmem_req_bits_size),
    .io_dmem_req_bits_signed(core_io_dmem_req_bits_signed),
    .io_dmem_s1_kill(core_io_dmem_s1_kill),
    .io_dmem_s1_data_data(core_io_dmem_s1_data_data),
    .io_dmem_s2_nack(core_io_dmem_s2_nack),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_size(core_io_dmem_resp_bits_size),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),
    .io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
    .io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),
    .io_dmem_replay_next(core_io_dmem_replay_next),
    .io_dmem_s2_xcpt_ma_ld(core_io_dmem_s2_xcpt_ma_ld),
    .io_dmem_s2_xcpt_ma_st(core_io_dmem_s2_xcpt_ma_st),
    .io_dmem_s2_xcpt_pf_ld(core_io_dmem_s2_xcpt_pf_ld),
    .io_dmem_s2_xcpt_pf_st(core_io_dmem_s2_xcpt_pf_st),
    .io_dmem_s2_xcpt_ae_ld(core_io_dmem_s2_xcpt_ae_ld),
    .io_dmem_s2_xcpt_ae_st(core_io_dmem_s2_xcpt_ae_st),
    .io_dmem_ordered(core_io_dmem_ordered),
    .io_dmem_perf_release(core_io_dmem_perf_release),
    .io_dmem_perf_grant(core_io_dmem_perf_grant),
    .io_ptw_ptbr_mode(core_io_ptw_ptbr_mode),
    .io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),
    .io_ptw_sfence_valid(core_io_ptw_sfence_valid),
    .io_ptw_sfence_bits_rs1(core_io_ptw_sfence_bits_rs1),
    .io_ptw_status_debug(core_io_ptw_status_debug),
    .io_ptw_status_dprv(core_io_ptw_status_dprv),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_mxr(core_io_ptw_status_mxr),
    .io_ptw_status_sum(core_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(core_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(core_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(core_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(core_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(core_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(core_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(core_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(core_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(core_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(core_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(core_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(core_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(core_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(core_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(core_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(core_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(core_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(core_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(core_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(core_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(core_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(core_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(core_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(core_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(core_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(core_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(core_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(core_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(core_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(core_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(core_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(core_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(core_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(core_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(core_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(core_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(core_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(core_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(core_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(core_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(core_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(core_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(core_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(core_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(core_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(core_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(core_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(core_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(core_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(core_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(core_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(core_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(core_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(core_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(core_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(core_io_ptw_pmp_7_mask),
    .io_ptw_customCSRs_csrs_0_value(core_io_ptw_customCSRs_csrs_0_value),
    .io_fpu_inst(core_io_fpu_inst),
    .io_fpu_fromint_data(core_io_fpu_fromint_data),
    .io_fpu_fcsr_rm(core_io_fpu_fcsr_rm),
    .io_fpu_fcsr_flags_valid(core_io_fpu_fcsr_flags_valid),
    .io_fpu_fcsr_flags_bits(core_io_fpu_fcsr_flags_bits),
    .io_fpu_store_data(core_io_fpu_store_data),
    .io_fpu_toint_data(core_io_fpu_toint_data),
    .io_fpu_dmem_resp_val(core_io_fpu_dmem_resp_val),
    .io_fpu_dmem_resp_type(core_io_fpu_dmem_resp_type),
    .io_fpu_dmem_resp_tag(core_io_fpu_dmem_resp_tag),
    .io_fpu_dmem_resp_data(core_io_fpu_dmem_resp_data),
    .io_fpu_valid(core_io_fpu_valid),
    .io_fpu_fcsr_rdy(core_io_fpu_fcsr_rdy),
    .io_fpu_nack_mem(core_io_fpu_nack_mem),
    .io_fpu_illegal_rm(core_io_fpu_illegal_rm),
    .io_fpu_killx(core_io_fpu_killx),
    .io_fpu_killm(core_io_fpu_killm),
    .io_fpu_dec_wen(core_io_fpu_dec_wen),
    .io_fpu_dec_ren1(core_io_fpu_dec_ren1),
    .io_fpu_dec_ren2(core_io_fpu_dec_ren2),
    .io_fpu_dec_ren3(core_io_fpu_dec_ren3),
    .io_fpu_sboard_set(core_io_fpu_sboard_set),
    .io_fpu_sboard_clr(core_io_fpu_sboard_clr),
    .io_fpu_sboard_clra(core_io_fpu_sboard_clra),
    .io_wfi(core_io_wfi),
    .io_covSum(core_io_covSum),
    .metaAssert(core_metaAssert),
    .metaReset(core_metaReset),
    .csr_halt(core_csr_halt),
    .div_halt(core_div_halt),
    .ibuf_halt(core_ibuf_halt),
    .Checking_Rocket_regstate(Rocket_regstate),		//Jaewon_Rocket_regstate
    .Checking_Rocket_covSum(Rocket_covSum)		//Jaewon_Rocket_regstat
  );
  assign auto_tl_master_xing_out_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_a_bits_param = buffer_auto_out_a_bits_param; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_a_bits_corrupt = buffer_auto_out_a_bits_corrupt; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_b_ready = buffer_auto_out_b_ready; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_c_valid = buffer_auto_out_c_valid; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_c_bits_opcode = buffer_auto_out_c_bits_opcode; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_c_bits_param = buffer_auto_out_c_bits_param; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_c_bits_size = buffer_auto_out_c_bits_size; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_c_bits_source = buffer_auto_out_c_bits_source; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_c_bits_address = buffer_auto_out_c_bits_address; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_c_bits_data = buffer_auto_out_c_bits_data; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_c_bits_corrupt = buffer_auto_out_c_bits_corrupt; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_e_valid = buffer_auto_out_e_valid; // @[LazyModule.scala 305:12]
  assign auto_tl_master_xing_out_e_bits_sink = buffer_auto_out_e_bits_sink; // @[LazyModule.scala 305:12]
  assign auto_wfi_out_0 = _T_33; // @[LazyModule.scala 305:12]
  assign auto_cease_out_0 = 1'h0; // @[LazyModule.scala 305:12]
  assign auto_halt_out_0 = 1'h0; // @[LazyModule.scala 305:12]
  assign tlMasterXbar_clock = clock;
  assign tlMasterXbar_reset = reset;
  assign tlMasterXbar_auto_in_1_a_valid = frontend_auto_icache_master_out_a_valid; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_1_a_bits_address = frontend_auto_icache_master_out_a_bits_address; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_a_valid = dcache_auto_out_a_valid; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_a_bits_opcode = dcache_auto_out_a_bits_opcode; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_a_bits_param = dcache_auto_out_a_bits_param; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_a_bits_size = dcache_auto_out_a_bits_size; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_a_bits_source = dcache_auto_out_a_bits_source; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_a_bits_address = dcache_auto_out_a_bits_address; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_a_bits_mask = dcache_auto_out_a_bits_mask; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_a_bits_data = dcache_auto_out_a_bits_data; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_b_ready = dcache_auto_out_b_ready; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_c_valid = dcache_auto_out_c_valid; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_c_bits_opcode = dcache_auto_out_c_bits_opcode; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_c_bits_param = dcache_auto_out_c_bits_param; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_c_bits_size = dcache_auto_out_c_bits_size; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_c_bits_source = dcache_auto_out_c_bits_source; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_c_bits_address = dcache_auto_out_c_bits_address; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_c_bits_data = dcache_auto_out_c_bits_data; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_d_ready = dcache_auto_out_d_ready; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_e_valid = dcache_auto_out_e_valid; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_in_0_e_bits_sink = dcache_auto_out_e_bits_sink; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_b_valid = buffer_auto_in_b_valid; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_b_bits_opcode = buffer_auto_in_b_bits_opcode; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_b_bits_param = buffer_auto_in_b_bits_param; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_b_bits_size = buffer_auto_in_b_bits_size; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_b_bits_source = buffer_auto_in_b_bits_source; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_b_bits_address = buffer_auto_in_b_bits_address; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_b_bits_mask = buffer_auto_in_b_bits_mask; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_b_bits_corrupt = buffer_auto_in_b_bits_corrupt; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_c_ready = buffer_auto_in_c_ready; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_d_bits_param = buffer_auto_in_d_bits_param; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 290:16]
  assign tlMasterXbar_auto_out_e_ready = buffer_auto_in_e_ready; // @[LazyModule.scala 290:16]
  assign intXbar_auto_int_in_3_0 = intsink_3_auto_out_0; // @[LazyModule.scala 292:16]
  assign intXbar_auto_int_in_2_0 = intsink_2_auto_out_0; // @[LazyModule.scala 292:16]
  assign intXbar_auto_int_in_1_0 = intsink_1_auto_out_0; // @[LazyModule.scala 292:16]
  assign intXbar_auto_int_in_1_1 = intsink_1_auto_out_1; // @[LazyModule.scala 292:16]
  assign intXbar_auto_int_in_0_0 = intsink_auto_out_0; // @[LazyModule.scala 292:16]
  assign hartIdNode_auto_in = auto_hartid_in; // @[LazyModule.scala 292:16]
  assign resetVectorNode_auto_in = auto_reset_vector_in; // @[LazyModule.scala 292:16]
  assign dcache_gated_clock = clock;
  assign dcache_reset = reset;
  assign dcache_auto_out_a_ready = tlMasterXbar_auto_in_0_a_ready; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_b_valid = tlMasterXbar_auto_in_0_b_valid; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_b_bits_param = tlMasterXbar_auto_in_0_b_bits_param; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_b_bits_size = tlMasterXbar_auto_in_0_b_bits_size; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_b_bits_source = tlMasterXbar_auto_in_0_b_bits_source; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_b_bits_address = tlMasterXbar_auto_in_0_b_bits_address; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_c_ready = tlMasterXbar_auto_in_0_c_ready; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_d_valid = tlMasterXbar_auto_in_0_d_valid; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_d_bits_opcode = tlMasterXbar_auto_in_0_d_bits_opcode; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_d_bits_param = tlMasterXbar_auto_in_0_d_bits_param; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_d_bits_size = tlMasterXbar_auto_in_0_d_bits_size; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_d_bits_source = tlMasterXbar_auto_in_0_d_bits_source; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_d_bits_sink = tlMasterXbar_auto_in_0_d_bits_sink; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_d_bits_denied = tlMasterXbar_auto_in_0_d_bits_denied; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_d_bits_data = tlMasterXbar_auto_in_0_d_bits_data; // @[LazyModule.scala 290:16]
  assign dcache_auto_out_e_ready = tlMasterXbar_auto_in_0_e_ready; // @[LazyModule.scala 290:16]
  assign dcache_io_cpu_req_valid = dcacheArb_io_mem_req_valid; // @[HellaCache.scala 265:30]
  assign dcache_io_cpu_req_bits_addr = dcacheArb_io_mem_req_bits_addr; // @[HellaCache.scala 265:30]
  assign dcache_io_cpu_req_bits_tag = dcacheArb_io_mem_req_bits_tag; // @[HellaCache.scala 265:30]
  assign dcache_io_cpu_req_bits_cmd = dcacheArb_io_mem_req_bits_cmd; // @[HellaCache.scala 265:30]
  assign dcache_io_cpu_req_bits_size = dcacheArb_io_mem_req_bits_size; // @[HellaCache.scala 265:30]
  assign dcache_io_cpu_req_bits_signed = dcacheArb_io_mem_req_bits_signed; // @[HellaCache.scala 265:30]
  assign dcache_io_cpu_req_bits_phys = dcacheArb_io_mem_req_bits_phys; // @[HellaCache.scala 265:30]
  assign dcache_io_cpu_s1_kill = dcacheArb_io_mem_s1_kill; // @[HellaCache.scala 265:30]
  assign dcache_io_cpu_s1_data_data = dcacheArb_io_mem_s1_data_data; // @[HellaCache.scala 265:30]
  assign dcache_io_ptw_req_ready = ptw_io_requestor_0_req_ready; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_valid = ptw_io_requestor_0_resp_valid; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_bits_ae = ptw_io_requestor_0_resp_bits_ae; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_bits_pte_ppn = ptw_io_requestor_0_resp_bits_pte_ppn; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_bits_pte_d = ptw_io_requestor_0_resp_bits_pte_d; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_bits_pte_a = ptw_io_requestor_0_resp_bits_pte_a; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_bits_pte_g = ptw_io_requestor_0_resp_bits_pte_g; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_bits_pte_u = ptw_io_requestor_0_resp_bits_pte_u; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_bits_pte_x = ptw_io_requestor_0_resp_bits_pte_x; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_bits_pte_w = ptw_io_requestor_0_resp_bits_pte_w; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_bits_pte_r = ptw_io_requestor_0_resp_bits_pte_r; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_bits_pte_v = ptw_io_requestor_0_resp_bits_pte_v; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_bits_level = ptw_io_requestor_0_resp_bits_level; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_resp_bits_homogeneous = ptw_io_requestor_0_resp_bits_homogeneous; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_ptbr_mode = ptw_io_requestor_0_ptbr_mode; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_status_debug = ptw_io_requestor_0_status_debug; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_status_dprv = ptw_io_requestor_0_status_dprv; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_status_mxr = ptw_io_requestor_0_status_mxr; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_status_sum = ptw_io_requestor_0_status_sum; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_0_cfg_l = ptw_io_requestor_0_pmp_0_cfg_l; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_0_cfg_a = ptw_io_requestor_0_pmp_0_cfg_a; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_0_cfg_x = ptw_io_requestor_0_pmp_0_cfg_x; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_0_cfg_w = ptw_io_requestor_0_pmp_0_cfg_w; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_0_cfg_r = ptw_io_requestor_0_pmp_0_cfg_r; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_0_addr = ptw_io_requestor_0_pmp_0_addr; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_0_mask = ptw_io_requestor_0_pmp_0_mask; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_1_cfg_l = ptw_io_requestor_0_pmp_1_cfg_l; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_1_cfg_a = ptw_io_requestor_0_pmp_1_cfg_a; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_1_cfg_x = ptw_io_requestor_0_pmp_1_cfg_x; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_1_cfg_w = ptw_io_requestor_0_pmp_1_cfg_w; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_1_cfg_r = ptw_io_requestor_0_pmp_1_cfg_r; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_1_addr = ptw_io_requestor_0_pmp_1_addr; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_1_mask = ptw_io_requestor_0_pmp_1_mask; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_2_cfg_l = ptw_io_requestor_0_pmp_2_cfg_l; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_2_cfg_a = ptw_io_requestor_0_pmp_2_cfg_a; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_2_cfg_x = ptw_io_requestor_0_pmp_2_cfg_x; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_2_cfg_w = ptw_io_requestor_0_pmp_2_cfg_w; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_2_cfg_r = ptw_io_requestor_0_pmp_2_cfg_r; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_2_addr = ptw_io_requestor_0_pmp_2_addr; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_2_mask = ptw_io_requestor_0_pmp_2_mask; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_3_cfg_l = ptw_io_requestor_0_pmp_3_cfg_l; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_3_cfg_a = ptw_io_requestor_0_pmp_3_cfg_a; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_3_cfg_x = ptw_io_requestor_0_pmp_3_cfg_x; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_3_cfg_w = ptw_io_requestor_0_pmp_3_cfg_w; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_3_cfg_r = ptw_io_requestor_0_pmp_3_cfg_r; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_3_addr = ptw_io_requestor_0_pmp_3_addr; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_3_mask = ptw_io_requestor_0_pmp_3_mask; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_4_cfg_l = ptw_io_requestor_0_pmp_4_cfg_l; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_4_cfg_a = ptw_io_requestor_0_pmp_4_cfg_a; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_4_cfg_x = ptw_io_requestor_0_pmp_4_cfg_x; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_4_cfg_w = ptw_io_requestor_0_pmp_4_cfg_w; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_4_cfg_r = ptw_io_requestor_0_pmp_4_cfg_r; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_4_addr = ptw_io_requestor_0_pmp_4_addr; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_4_mask = ptw_io_requestor_0_pmp_4_mask; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_5_cfg_l = ptw_io_requestor_0_pmp_5_cfg_l; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_5_cfg_a = ptw_io_requestor_0_pmp_5_cfg_a; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_5_cfg_x = ptw_io_requestor_0_pmp_5_cfg_x; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_5_cfg_w = ptw_io_requestor_0_pmp_5_cfg_w; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_5_cfg_r = ptw_io_requestor_0_pmp_5_cfg_r; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_5_addr = ptw_io_requestor_0_pmp_5_addr; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_5_mask = ptw_io_requestor_0_pmp_5_mask; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_6_cfg_l = ptw_io_requestor_0_pmp_6_cfg_l; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_6_cfg_a = ptw_io_requestor_0_pmp_6_cfg_a; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_6_cfg_x = ptw_io_requestor_0_pmp_6_cfg_x; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_6_cfg_w = ptw_io_requestor_0_pmp_6_cfg_w; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_6_cfg_r = ptw_io_requestor_0_pmp_6_cfg_r; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_6_addr = ptw_io_requestor_0_pmp_6_addr; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_6_mask = ptw_io_requestor_0_pmp_6_mask; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_7_cfg_l = ptw_io_requestor_0_pmp_7_cfg_l; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_7_cfg_a = ptw_io_requestor_0_pmp_7_cfg_a; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_7_cfg_x = ptw_io_requestor_0_pmp_7_cfg_x; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_7_cfg_w = ptw_io_requestor_0_pmp_7_cfg_w; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_7_cfg_r = ptw_io_requestor_0_pmp_7_cfg_r; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_7_addr = ptw_io_requestor_0_pmp_7_addr; // @[RocketTile.scala 191:20]
  assign dcache_io_ptw_pmp_7_mask = ptw_io_requestor_0_pmp_7_mask; // @[RocketTile.scala 191:20]
  assign frontend_gated_clock = clock;
  assign frontend_reset = reset;
  assign frontend_auto_icache_master_out_a_ready = tlMasterXbar_auto_in_1_a_ready; // @[LazyModule.scala 290:16]
  assign frontend_auto_icache_master_out_d_valid = tlMasterXbar_auto_in_1_d_valid; // @[LazyModule.scala 290:16]
  assign frontend_auto_icache_master_out_d_bits_opcode = tlMasterXbar_auto_in_1_d_bits_opcode; // @[LazyModule.scala 290:16]
  assign frontend_auto_icache_master_out_d_bits_size = tlMasterXbar_auto_in_1_d_bits_size; // @[LazyModule.scala 290:16]
  assign frontend_auto_icache_master_out_d_bits_data = tlMasterXbar_auto_in_1_d_bits_data; // @[LazyModule.scala 290:16]
  assign frontend_auto_icache_master_out_d_bits_corrupt = tlMasterXbar_auto_in_1_d_bits_corrupt; // @[LazyModule.scala 290:16]
  assign frontend_auto_reset_vector_sink_in = resetVectorNode_auto_out_1; // @[LazyModule.scala 292:16]
  assign frontend_io_cpu_might_request = core_io_imem_might_request; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_req_valid = core_io_imem_req_valid; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_req_bits_pc = core_io_imem_req_bits_pc; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_req_bits_speculative = core_io_imem_req_bits_speculative; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_sfence_valid = core_io_imem_sfence_valid; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_sfence_bits_rs1 = core_io_imem_sfence_bits_rs1; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_sfence_bits_rs2 = core_io_imem_sfence_bits_rs2; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_sfence_bits_addr = core_io_imem_sfence_bits_addr; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_resp_ready = core_io_imem_resp_ready; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_btb_update_valid = core_io_imem_btb_update_valid; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_btb_update_bits_prediction_entry = core_io_imem_btb_update_bits_prediction_entry; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_btb_update_bits_pc = core_io_imem_btb_update_bits_pc; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_btb_update_bits_isValid = core_io_imem_btb_update_bits_isValid; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_btb_update_bits_br_pc = core_io_imem_btb_update_bits_br_pc; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_btb_update_bits_cfiType = core_io_imem_btb_update_bits_cfiType; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_bht_update_valid = core_io_imem_bht_update_valid; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_bht_update_bits_prediction_history = core_io_imem_bht_update_bits_prediction_history; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_bht_update_bits_pc = core_io_imem_bht_update_bits_pc; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_bht_update_bits_branch = core_io_imem_bht_update_bits_branch; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_bht_update_bits_taken = core_io_imem_bht_update_bits_taken; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_bht_update_bits_mispredict = core_io_imem_bht_update_bits_mispredict; // @[RocketTile.scala 166:32]
  assign frontend_io_cpu_flush_icache = core_io_imem_flush_icache; // @[RocketTile.scala 166:32]
  assign frontend_io_ptw_req_ready = ptw_io_requestor_1_req_ready; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_valid = ptw_io_requestor_1_resp_valid; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_bits_ae = ptw_io_requestor_1_resp_bits_ae; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_bits_pte_ppn = ptw_io_requestor_1_resp_bits_pte_ppn; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_bits_pte_d = ptw_io_requestor_1_resp_bits_pte_d; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_bits_pte_a = ptw_io_requestor_1_resp_bits_pte_a; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_bits_pte_g = ptw_io_requestor_1_resp_bits_pte_g; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_bits_pte_u = ptw_io_requestor_1_resp_bits_pte_u; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_bits_pte_x = ptw_io_requestor_1_resp_bits_pte_x; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_bits_pte_w = ptw_io_requestor_1_resp_bits_pte_w; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_bits_pte_r = ptw_io_requestor_1_resp_bits_pte_r; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_bits_pte_v = ptw_io_requestor_1_resp_bits_pte_v; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_bits_level = ptw_io_requestor_1_resp_bits_level; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_resp_bits_homogeneous = ptw_io_requestor_1_resp_bits_homogeneous; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_ptbr_mode = ptw_io_requestor_1_ptbr_mode; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_status_debug = ptw_io_requestor_1_status_debug; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_status_prv = ptw_io_requestor_1_status_prv; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_0_cfg_l = ptw_io_requestor_1_pmp_0_cfg_l; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_0_cfg_a = ptw_io_requestor_1_pmp_0_cfg_a; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_0_cfg_x = ptw_io_requestor_1_pmp_0_cfg_x; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_0_cfg_w = ptw_io_requestor_1_pmp_0_cfg_w; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_0_cfg_r = ptw_io_requestor_1_pmp_0_cfg_r; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_0_addr = ptw_io_requestor_1_pmp_0_addr; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_0_mask = ptw_io_requestor_1_pmp_0_mask; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_1_cfg_l = ptw_io_requestor_1_pmp_1_cfg_l; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_1_cfg_a = ptw_io_requestor_1_pmp_1_cfg_a; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_1_cfg_x = ptw_io_requestor_1_pmp_1_cfg_x; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_1_cfg_w = ptw_io_requestor_1_pmp_1_cfg_w; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_1_cfg_r = ptw_io_requestor_1_pmp_1_cfg_r; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_1_addr = ptw_io_requestor_1_pmp_1_addr; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_1_mask = ptw_io_requestor_1_pmp_1_mask; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_2_cfg_l = ptw_io_requestor_1_pmp_2_cfg_l; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_2_cfg_a = ptw_io_requestor_1_pmp_2_cfg_a; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_2_cfg_x = ptw_io_requestor_1_pmp_2_cfg_x; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_2_cfg_w = ptw_io_requestor_1_pmp_2_cfg_w; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_2_cfg_r = ptw_io_requestor_1_pmp_2_cfg_r; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_2_addr = ptw_io_requestor_1_pmp_2_addr; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_2_mask = ptw_io_requestor_1_pmp_2_mask; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_3_cfg_l = ptw_io_requestor_1_pmp_3_cfg_l; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_3_cfg_a = ptw_io_requestor_1_pmp_3_cfg_a; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_3_cfg_x = ptw_io_requestor_1_pmp_3_cfg_x; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_3_cfg_w = ptw_io_requestor_1_pmp_3_cfg_w; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_3_cfg_r = ptw_io_requestor_1_pmp_3_cfg_r; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_3_addr = ptw_io_requestor_1_pmp_3_addr; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_3_mask = ptw_io_requestor_1_pmp_3_mask; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_4_cfg_l = ptw_io_requestor_1_pmp_4_cfg_l; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_4_cfg_a = ptw_io_requestor_1_pmp_4_cfg_a; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_4_cfg_x = ptw_io_requestor_1_pmp_4_cfg_x; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_4_cfg_w = ptw_io_requestor_1_pmp_4_cfg_w; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_4_cfg_r = ptw_io_requestor_1_pmp_4_cfg_r; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_4_addr = ptw_io_requestor_1_pmp_4_addr; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_4_mask = ptw_io_requestor_1_pmp_4_mask; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_5_cfg_l = ptw_io_requestor_1_pmp_5_cfg_l; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_5_cfg_a = ptw_io_requestor_1_pmp_5_cfg_a; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_5_cfg_x = ptw_io_requestor_1_pmp_5_cfg_x; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_5_cfg_w = ptw_io_requestor_1_pmp_5_cfg_w; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_5_cfg_r = ptw_io_requestor_1_pmp_5_cfg_r; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_5_addr = ptw_io_requestor_1_pmp_5_addr; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_5_mask = ptw_io_requestor_1_pmp_5_mask; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_6_cfg_l = ptw_io_requestor_1_pmp_6_cfg_l; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_6_cfg_a = ptw_io_requestor_1_pmp_6_cfg_a; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_6_cfg_x = ptw_io_requestor_1_pmp_6_cfg_x; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_6_cfg_w = ptw_io_requestor_1_pmp_6_cfg_w; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_6_cfg_r = ptw_io_requestor_1_pmp_6_cfg_r; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_6_addr = ptw_io_requestor_1_pmp_6_addr; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_6_mask = ptw_io_requestor_1_pmp_6_mask; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_7_cfg_l = ptw_io_requestor_1_pmp_7_cfg_l; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_7_cfg_a = ptw_io_requestor_1_pmp_7_cfg_a; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_7_cfg_x = ptw_io_requestor_1_pmp_7_cfg_x; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_7_cfg_w = ptw_io_requestor_1_pmp_7_cfg_w; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_7_cfg_r = ptw_io_requestor_1_pmp_7_cfg_r; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_7_addr = ptw_io_requestor_1_pmp_7_addr; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_pmp_7_mask = ptw_io_requestor_1_pmp_7_mask; // @[RocketTile.scala 191:20]
  assign frontend_io_ptw_customCSRs_csrs_0_value = ptw_io_requestor_1_customCSRs_csrs_0_value; // @[RocketTile.scala 191:20]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_auto_in_a_valid = tlMasterXbar_auto_out_a_valid; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_a_bits_opcode = tlMasterXbar_auto_out_a_bits_opcode; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_a_bits_param = tlMasterXbar_auto_out_a_bits_param; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_a_bits_size = tlMasterXbar_auto_out_a_bits_size; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_a_bits_source = tlMasterXbar_auto_out_a_bits_source; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_a_bits_address = tlMasterXbar_auto_out_a_bits_address; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_a_bits_mask = tlMasterXbar_auto_out_a_bits_mask; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_a_bits_data = tlMasterXbar_auto_out_a_bits_data; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_a_bits_corrupt = tlMasterXbar_auto_out_a_bits_corrupt; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_b_ready = tlMasterXbar_auto_out_b_ready; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_c_valid = tlMasterXbar_auto_out_c_valid; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_c_bits_opcode = tlMasterXbar_auto_out_c_bits_opcode; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_c_bits_param = tlMasterXbar_auto_out_c_bits_param; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_c_bits_size = tlMasterXbar_auto_out_c_bits_size; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_c_bits_source = tlMasterXbar_auto_out_c_bits_source; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_c_bits_address = tlMasterXbar_auto_out_c_bits_address; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_c_bits_data = tlMasterXbar_auto_out_c_bits_data; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_d_ready = tlMasterXbar_auto_out_d_ready; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_e_valid = tlMasterXbar_auto_out_e_valid; // @[LazyModule.scala 292:16]
  assign buffer_auto_in_e_bits_sink = tlMasterXbar_auto_out_e_bits_sink; // @[LazyModule.scala 292:16]
  assign buffer_auto_out_a_ready = auto_tl_master_xing_out_a_ready; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_b_valid = auto_tl_master_xing_out_b_valid; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_b_bits_opcode = auto_tl_master_xing_out_b_bits_opcode; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_b_bits_param = auto_tl_master_xing_out_b_bits_param; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_b_bits_size = auto_tl_master_xing_out_b_bits_size; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_b_bits_source = auto_tl_master_xing_out_b_bits_source; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_b_bits_address = auto_tl_master_xing_out_b_bits_address; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_b_bits_mask = auto_tl_master_xing_out_b_bits_mask; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_b_bits_corrupt = auto_tl_master_xing_out_b_bits_corrupt; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_c_ready = auto_tl_master_xing_out_c_ready; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_d_valid = auto_tl_master_xing_out_d_valid; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_d_bits_opcode = auto_tl_master_xing_out_d_bits_opcode; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_d_bits_param = auto_tl_master_xing_out_d_bits_param; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_d_bits_size = auto_tl_master_xing_out_d_bits_size; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_d_bits_source = auto_tl_master_xing_out_d_bits_source; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_d_bits_sink = auto_tl_master_xing_out_d_bits_sink; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_d_bits_denied = auto_tl_master_xing_out_d_bits_denied; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_d_bits_data = auto_tl_master_xing_out_d_bits_data; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_d_bits_corrupt = auto_tl_master_xing_out_d_bits_corrupt; // @[LazyModule.scala 290:16]
  assign buffer_auto_out_e_ready = auto_tl_master_xing_out_e_ready; // @[LazyModule.scala 290:16]
  assign intsink_clock = clock;
  assign intsink_auto_in_sync_0 = auto_intsink_in_sync_0; // @[LazyModule.scala 303:16]
  assign intsink_1_auto_in_sync_0 = auto_int_in_xing_in_0_sync_0; // @[LazyModule.scala 292:16]
  assign intsink_1_auto_in_sync_1 = auto_int_in_xing_in_0_sync_1; // @[LazyModule.scala 292:16]
  assign intsink_2_auto_in_sync_0 = auto_int_in_xing_in_1_sync_0; // @[LazyModule.scala 292:16]
  assign intsink_3_auto_in_sync_0 = auto_int_in_xing_in_2_sync_0; // @[LazyModule.scala 292:16]
  assign fpuOpt_clock = clock;
  assign fpuOpt_reset = reset;
  assign fpuOpt_io_inst = core_io_fpu_inst; // @[RocketTile.scala 168:39]
  assign fpuOpt_io_fromint_data = core_io_fpu_fromint_data; // @[RocketTile.scala 168:39]
  assign fpuOpt_io_fcsr_rm = core_io_fpu_fcsr_rm; // @[RocketTile.scala 168:39]
  assign fpuOpt_io_dmem_resp_val = core_io_fpu_dmem_resp_val; // @[RocketTile.scala 168:39]
  assign fpuOpt_io_dmem_resp_type = core_io_fpu_dmem_resp_type; // @[RocketTile.scala 168:39]
  assign fpuOpt_io_dmem_resp_tag = core_io_fpu_dmem_resp_tag; // @[RocketTile.scala 168:39]
  assign fpuOpt_io_dmem_resp_data = core_io_fpu_dmem_resp_data; // @[RocketTile.scala 168:39]
  assign fpuOpt_io_valid = core_io_fpu_valid; // @[RocketTile.scala 168:39]
  assign fpuOpt_io_killx = core_io_fpu_killx; // @[RocketTile.scala 168:39]
  assign fpuOpt_io_killm = core_io_fpu_killm; // @[RocketTile.scala 168:39]
  assign dcacheArb_clock = clock;
  assign dcacheArb_io_requestor_0_req_valid = ptw_io_mem_req_valid; // @[RocketTile.scala 190:26]
  assign dcacheArb_io_requestor_0_req_bits_addr = ptw_io_mem_req_bits_addr; // @[RocketTile.scala 190:26]
  assign dcacheArb_io_requestor_0_s1_kill = ptw_io_mem_s1_kill; // @[RocketTile.scala 190:26]
  assign dcacheArb_io_requestor_1_req_valid = core_io_dmem_req_valid; // @[RocketTile.scala 190:26]
  assign dcacheArb_io_requestor_1_req_bits_addr = core_io_dmem_req_bits_addr; // @[RocketTile.scala 190:26]
  assign dcacheArb_io_requestor_1_req_bits_tag = core_io_dmem_req_bits_tag; // @[RocketTile.scala 190:26]
  assign dcacheArb_io_requestor_1_req_bits_cmd = core_io_dmem_req_bits_cmd; // @[RocketTile.scala 190:26]
  assign dcacheArb_io_requestor_1_req_bits_size = core_io_dmem_req_bits_size; // @[RocketTile.scala 190:26]
  assign dcacheArb_io_requestor_1_req_bits_signed = core_io_dmem_req_bits_signed; // @[RocketTile.scala 190:26]
  assign dcacheArb_io_requestor_1_s1_kill = core_io_dmem_s1_kill; // @[RocketTile.scala 190:26]
  assign dcacheArb_io_requestor_1_s1_data_data = core_io_dmem_s1_data_data; // @[RocketTile.scala 190:26]
  assign dcacheArb_io_mem_req_ready = dcache_io_cpu_req_ready; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_s2_nack = dcache_io_cpu_s2_nack; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_resp_valid = dcache_io_cpu_resp_valid; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_resp_bits_tag = dcache_io_cpu_resp_bits_tag; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_resp_bits_size = dcache_io_cpu_resp_bits_size; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_resp_bits_data = dcache_io_cpu_resp_bits_data; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_resp_bits_replay = dcache_io_cpu_resp_bits_replay; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_resp_bits_has_data = dcache_io_cpu_resp_bits_has_data; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_resp_bits_data_word_bypass = dcache_io_cpu_resp_bits_data_word_bypass; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_replay_next = dcache_io_cpu_replay_next; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_s2_xcpt_ma_ld = dcache_io_cpu_s2_xcpt_ma_ld; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_s2_xcpt_ma_st = dcache_io_cpu_s2_xcpt_ma_st; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_s2_xcpt_pf_ld = dcache_io_cpu_s2_xcpt_pf_ld; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_s2_xcpt_pf_st = dcache_io_cpu_s2_xcpt_pf_st; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_s2_xcpt_ae_ld = dcache_io_cpu_s2_xcpt_ae_ld; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_s2_xcpt_ae_st = dcache_io_cpu_s2_xcpt_ae_st; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_ordered = dcache_io_cpu_ordered; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_perf_release = dcache_io_cpu_perf_release; // @[HellaCache.scala 265:30]
  assign dcacheArb_io_mem_perf_grant = dcache_io_cpu_perf_grant; // @[HellaCache.scala 265:30]
  assign ptw_clock = clock;
  assign ptw_reset = reset;
  assign ptw_io_requestor_0_req_valid = dcache_io_ptw_req_valid; // @[RocketTile.scala 191:20]
  assign ptw_io_requestor_0_req_bits_bits_addr = dcache_io_ptw_req_bits_bits_addr; // @[RocketTile.scala 191:20]
  assign ptw_io_requestor_1_req_valid = frontend_io_ptw_req_valid; // @[RocketTile.scala 191:20]
  assign ptw_io_requestor_1_req_bits_valid = frontend_io_ptw_req_bits_valid; // @[RocketTile.scala 191:20]
  assign ptw_io_requestor_1_req_bits_bits_addr = frontend_io_ptw_req_bits_bits_addr; // @[RocketTile.scala 191:20]
  assign ptw_io_mem_req_ready = dcacheArb_io_requestor_0_req_ready; // @[RocketTile.scala 190:26]
  assign ptw_io_mem_s2_nack = dcacheArb_io_requestor_0_s2_nack; // @[RocketTile.scala 190:26]
  assign ptw_io_mem_resp_valid = dcacheArb_io_requestor_0_resp_valid; // @[RocketTile.scala 190:26]
  assign ptw_io_mem_resp_bits_data = dcacheArb_io_requestor_0_resp_bits_data; // @[RocketTile.scala 190:26]
  assign ptw_io_mem_s2_xcpt_ae_ld = dcacheArb_io_requestor_0_s2_xcpt_ae_ld; // @[RocketTile.scala 190:26]
  assign ptw_io_dpath_ptbr_mode = core_io_ptw_ptbr_mode; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_ptbr_ppn = core_io_ptw_ptbr_ppn; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_sfence_valid = core_io_ptw_sfence_valid; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_sfence_bits_rs1 = core_io_ptw_sfence_bits_rs1; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_status_debug = core_io_ptw_status_debug; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_status_dprv = core_io_ptw_status_dprv; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_status_prv = core_io_ptw_status_prv; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_status_mxr = core_io_ptw_status_mxr; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_status_sum = core_io_ptw_status_sum; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_0_cfg_l = core_io_ptw_pmp_0_cfg_l; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_0_cfg_a = core_io_ptw_pmp_0_cfg_a; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_0_cfg_x = core_io_ptw_pmp_0_cfg_x; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_0_cfg_w = core_io_ptw_pmp_0_cfg_w; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_0_cfg_r = core_io_ptw_pmp_0_cfg_r; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_0_addr = core_io_ptw_pmp_0_addr; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_0_mask = core_io_ptw_pmp_0_mask; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_1_cfg_l = core_io_ptw_pmp_1_cfg_l; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_1_cfg_a = core_io_ptw_pmp_1_cfg_a; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_1_cfg_x = core_io_ptw_pmp_1_cfg_x; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_1_cfg_w = core_io_ptw_pmp_1_cfg_w; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_1_cfg_r = core_io_ptw_pmp_1_cfg_r; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_1_addr = core_io_ptw_pmp_1_addr; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_1_mask = core_io_ptw_pmp_1_mask; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_2_cfg_l = core_io_ptw_pmp_2_cfg_l; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_2_cfg_a = core_io_ptw_pmp_2_cfg_a; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_2_cfg_x = core_io_ptw_pmp_2_cfg_x; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_2_cfg_w = core_io_ptw_pmp_2_cfg_w; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_2_cfg_r = core_io_ptw_pmp_2_cfg_r; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_2_addr = core_io_ptw_pmp_2_addr; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_2_mask = core_io_ptw_pmp_2_mask; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_3_cfg_l = core_io_ptw_pmp_3_cfg_l; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_3_cfg_a = core_io_ptw_pmp_3_cfg_a; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_3_cfg_x = core_io_ptw_pmp_3_cfg_x; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_3_cfg_w = core_io_ptw_pmp_3_cfg_w; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_3_cfg_r = core_io_ptw_pmp_3_cfg_r; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_3_addr = core_io_ptw_pmp_3_addr; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_3_mask = core_io_ptw_pmp_3_mask; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_4_cfg_l = core_io_ptw_pmp_4_cfg_l; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_4_cfg_a = core_io_ptw_pmp_4_cfg_a; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_4_cfg_x = core_io_ptw_pmp_4_cfg_x; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_4_cfg_w = core_io_ptw_pmp_4_cfg_w; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_4_cfg_r = core_io_ptw_pmp_4_cfg_r; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_4_addr = core_io_ptw_pmp_4_addr; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_4_mask = core_io_ptw_pmp_4_mask; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_5_cfg_l = core_io_ptw_pmp_5_cfg_l; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_5_cfg_a = core_io_ptw_pmp_5_cfg_a; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_5_cfg_x = core_io_ptw_pmp_5_cfg_x; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_5_cfg_w = core_io_ptw_pmp_5_cfg_w; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_5_cfg_r = core_io_ptw_pmp_5_cfg_r; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_5_addr = core_io_ptw_pmp_5_addr; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_5_mask = core_io_ptw_pmp_5_mask; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_6_cfg_l = core_io_ptw_pmp_6_cfg_l; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_6_cfg_a = core_io_ptw_pmp_6_cfg_a; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_6_cfg_x = core_io_ptw_pmp_6_cfg_x; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_6_cfg_w = core_io_ptw_pmp_6_cfg_w; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_6_cfg_r = core_io_ptw_pmp_6_cfg_r; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_6_addr = core_io_ptw_pmp_6_addr; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_6_mask = core_io_ptw_pmp_6_mask; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_7_cfg_l = core_io_ptw_pmp_7_cfg_l; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_7_cfg_a = core_io_ptw_pmp_7_cfg_a; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_7_cfg_x = core_io_ptw_pmp_7_cfg_x; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_7_cfg_w = core_io_ptw_pmp_7_cfg_w; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_7_cfg_r = core_io_ptw_pmp_7_cfg_r; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_7_addr = core_io_ptw_pmp_7_addr; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_pmp_7_mask = core_io_ptw_pmp_7_mask; // @[RocketTile.scala 169:15]
  assign ptw_io_dpath_customCSRs_csrs_0_value = core_io_ptw_customCSRs_csrs_0_value; // @[RocketTile.scala 169:15]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_hartid = hartIdNode_auto_out_0; // @[RocketTile.scala 161:18]
  assign core_io_interrupts_debug = intXbar_auto_int_out_0; // @[Interrupts.scala 75:93]
  assign core_io_interrupts_mtip = intXbar_auto_int_out_2; // @[Interrupts.scala 75:93]
  assign core_io_interrupts_msip = intXbar_auto_int_out_1; // @[Interrupts.scala 75:93]
  assign core_io_interrupts_meip = intXbar_auto_int_out_3; // @[Interrupts.scala 75:93]
  assign core_io_interrupts_seip = intXbar_auto_int_out_4; // @[Interrupts.scala 75:93]
  assign core_io_imem_resp_valid = frontend_io_cpu_resp_valid; // @[RocketTile.scala 166:32]
  assign core_io_imem_resp_bits_btb_taken = frontend_io_cpu_resp_bits_btb_taken; // @[RocketTile.scala 166:32]
  assign core_io_imem_resp_bits_btb_bridx = frontend_io_cpu_resp_bits_btb_bridx; // @[RocketTile.scala 166:32]
  assign core_io_imem_resp_bits_btb_entry = frontend_io_cpu_resp_bits_btb_entry; // @[RocketTile.scala 166:32]
  assign core_io_imem_resp_bits_btb_bht_history = frontend_io_cpu_resp_bits_btb_bht_history; // @[RocketTile.scala 166:32]
  assign core_io_imem_resp_bits_pc = frontend_io_cpu_resp_bits_pc; // @[RocketTile.scala 166:32]
  assign core_io_imem_resp_bits_data = frontend_io_cpu_resp_bits_data; // @[RocketTile.scala 166:32]
  assign core_io_imem_resp_bits_xcpt_pf_inst = frontend_io_cpu_resp_bits_xcpt_pf_inst; // @[RocketTile.scala 166:32]
  assign core_io_imem_resp_bits_xcpt_ae_inst = frontend_io_cpu_resp_bits_xcpt_ae_inst; // @[RocketTile.scala 166:32]
  assign core_io_imem_resp_bits_replay = frontend_io_cpu_resp_bits_replay; // @[RocketTile.scala 166:32]
  assign core_io_dmem_req_ready = dcacheArb_io_requestor_1_req_ready; // @[RocketTile.scala 190:26]
  assign core_io_dmem_s2_nack = dcacheArb_io_requestor_1_s2_nack; // @[RocketTile.scala 190:26]
  assign core_io_dmem_resp_valid = dcacheArb_io_requestor_1_resp_valid; // @[RocketTile.scala 190:26]
  assign core_io_dmem_resp_bits_tag = dcacheArb_io_requestor_1_resp_bits_tag; // @[RocketTile.scala 190:26]
  assign core_io_dmem_resp_bits_size = dcacheArb_io_requestor_1_resp_bits_size; // @[RocketTile.scala 190:26]
  assign core_io_dmem_resp_bits_data = dcacheArb_io_requestor_1_resp_bits_data; // @[RocketTile.scala 190:26]
  assign core_io_dmem_resp_bits_replay = dcacheArb_io_requestor_1_resp_bits_replay; // @[RocketTile.scala 190:26]
  assign core_io_dmem_resp_bits_has_data = dcacheArb_io_requestor_1_resp_bits_has_data; // @[RocketTile.scala 190:26]
  assign core_io_dmem_resp_bits_data_word_bypass = dcacheArb_io_requestor_1_resp_bits_data_word_bypass; // @[RocketTile.scala 190:26]
  assign core_io_dmem_replay_next = dcacheArb_io_requestor_1_replay_next; // @[RocketTile.scala 190:26]
  assign core_io_dmem_s2_xcpt_ma_ld = dcacheArb_io_requestor_1_s2_xcpt_ma_ld; // @[RocketTile.scala 190:26]
  assign core_io_dmem_s2_xcpt_ma_st = dcacheArb_io_requestor_1_s2_xcpt_ma_st; // @[RocketTile.scala 190:26]
  assign core_io_dmem_s2_xcpt_pf_ld = dcacheArb_io_requestor_1_s2_xcpt_pf_ld; // @[RocketTile.scala 190:26]
  assign core_io_dmem_s2_xcpt_pf_st = dcacheArb_io_requestor_1_s2_xcpt_pf_st; // @[RocketTile.scala 190:26]
  assign core_io_dmem_s2_xcpt_ae_ld = dcacheArb_io_requestor_1_s2_xcpt_ae_ld; // @[RocketTile.scala 190:26]
  assign core_io_dmem_s2_xcpt_ae_st = dcacheArb_io_requestor_1_s2_xcpt_ae_st; // @[RocketTile.scala 190:26]
  assign core_io_dmem_ordered = dcacheArb_io_requestor_1_ordered; // @[RocketTile.scala 190:26]
  assign core_io_dmem_perf_release = dcacheArb_io_requestor_1_perf_release; // @[RocketTile.scala 190:26]
  assign core_io_dmem_perf_grant = dcacheArb_io_requestor_1_perf_grant; // @[RocketTile.scala 190:26]
  assign core_io_fpu_fcsr_flags_valid = fpuOpt_io_fcsr_flags_valid; // @[RocketTile.scala 168:39]
  assign core_io_fpu_fcsr_flags_bits = fpuOpt_io_fcsr_flags_bits; // @[RocketTile.scala 168:39]
  assign core_io_fpu_store_data = fpuOpt_io_store_data; // @[RocketTile.scala 168:39]
  assign core_io_fpu_toint_data = fpuOpt_io_toint_data; // @[RocketTile.scala 168:39]
  assign core_io_fpu_fcsr_rdy = fpuOpt_io_fcsr_rdy; // @[RocketTile.scala 168:39]
  assign core_io_fpu_nack_mem = fpuOpt_io_nack_mem; // @[RocketTile.scala 168:39]
  assign core_io_fpu_illegal_rm = fpuOpt_io_illegal_rm; // @[RocketTile.scala 168:39]
  assign core_io_fpu_dec_wen = fpuOpt_io_dec_wen; // @[RocketTile.scala 168:39]
  assign core_io_fpu_dec_ren1 = fpuOpt_io_dec_ren1; // @[RocketTile.scala 168:39]
  assign core_io_fpu_dec_ren2 = fpuOpt_io_dec_ren2; // @[RocketTile.scala 168:39]
  assign core_io_fpu_dec_ren3 = fpuOpt_io_dec_ren3; // @[RocketTile.scala 168:39]
  assign core_io_fpu_sboard_set = fpuOpt_io_sboard_set; // @[RocketTile.scala 168:39]
  assign core_io_fpu_sboard_clr = fpuOpt_io_sboard_clr; // @[RocketTile.scala 168:39]
  assign core_io_fpu_sboard_clra = fpuOpt_io_sboard_clra; // @[RocketTile.scala 168:39]
  assign RocketTile_covSum = 30'h0;
  assign ptw_sum = RocketTile_covSum + ptw_io_covSum;
  assign resetVectorNode_sum = ptw_sum + resetVectorNode_io_covSum;
  assign dcacheArb_sum = resetVectorNode_sum + dcacheArb_io_covSum;
  assign tlMasterXbar_sum = dcacheArb_sum + tlMasterXbar_io_covSum;
  assign dcache_sum = tlMasterXbar_sum + dcache_io_covSum;
  assign intsink_3_sum = dcache_sum + intsink_3_io_covSum;
  assign intsink_1_sum = intsink_3_sum + intsink_1_io_covSum;
  assign buffer_sum = intsink_1_sum + buffer_io_covSum;
  assign core_sum = buffer_sum + core_io_covSum;
  assign fpuOpt_sum = core_sum + fpuOpt_io_covSum;
  assign intXbar_sum = fpuOpt_sum + intXbar_io_covSum;
  assign frontend_sum = intXbar_sum + frontend_io_covSum;
  assign hartIdNode_sum = frontend_sum + hartIdNode_io_covSum;
  assign intsink_sum = hartIdNode_sum + intsink_io_covSum;
  assign intsink_2_sum = intsink_sum + intsink_2_io_covSum;
  assign io_covSum = intsink_2_sum;
  assign intsink_1_metaAssert_wire = intsink_1_metaAssert;
  assign intsink_3_metaAssert_wire = intsink_3_metaAssert;
  assign intsink_metaAssert_wire = intsink_metaAssert;
  assign dcache_metaAssert_wire = dcache_metaAssert;
  assign intXbar_metaAssert_wire = intXbar_metaAssert;
  assign tlMasterXbar_metaAssert_wire = tlMasterXbar_metaAssert;
  assign frontend_metaAssert_wire = frontend_metaAssert;
  assign dcacheArb_metaAssert_wire = dcacheArb_metaAssert;
  assign buffer_metaAssert_wire = buffer_metaAssert;
  assign hartIdNode_metaAssert_wire = hartIdNode_metaAssert;
  assign fpuOpt_metaAssert_wire = fpuOpt_metaAssert;
  assign intsink_2_metaAssert_wire = intsink_2_metaAssert;
  assign resetVectorNode_metaAssert_wire = resetVectorNode_metaAssert;
  assign core_metaAssert_wire = core_metaAssert;
  assign ptw_metaAssert_wire = ptw_metaAssert;
  assign RocketTile_or8 = tlMasterXbar_metaAssert_wire | frontend_metaAssert_wire;
  assign RocketTile_or3 = hartIdNode_metaAssert_wire | RocketTile_or8;
  assign RocketTile_or9 = dcache_metaAssert_wire | fpuOpt_metaAssert_wire;
  assign RocketTile_or10 = intXbar_metaAssert_wire | ptw_metaAssert_wire;
  assign RocketTile_or4 = RocketTile_or9 | RocketTile_or10;
  assign RocketTile_or1 = RocketTile_or3 | RocketTile_or4;
  assign RocketTile_or11 = intsink_1_metaAssert_wire | intsink_2_metaAssert_wire;
  assign RocketTile_or12 = intsink_3_metaAssert_wire | core_metaAssert_wire;
  assign RocketTile_or5 = RocketTile_or11 | RocketTile_or12;
  assign RocketTile_or13 = dcacheArb_metaAssert_wire | intsink_metaAssert_wire;
  assign RocketTile_or14 = buffer_metaAssert_wire | resetVectorNode_metaAssert_wire;
  assign RocketTile_or6 = RocketTile_or13 | RocketTile_or14;
  assign RocketTile_or2 = RocketTile_or5 | RocketTile_or6;
  assign RocketTile_or0 = RocketTile_or1 | RocketTile_or2;
  assign metaAssert = RocketTile_metaAssert;
  assign ptw_metaReset = metaReset | ptw_halt;
  assign dcacheArb_metaReset = metaReset | dcacheArb_halt;
  assign tlMasterXbar_metaReset = metaReset | tlMasterXbar_halt;
  assign dcache_metaReset = metaReset | dcache_halt;
  assign buffer_metaReset = metaReset | buffer_halt;
  assign core_metaReset = metaReset | core_halt;
  assign fpuOpt_metaReset = metaReset | fpuOpt_halt;
  assign frontend_metaReset = metaReset | frontend_halt;
  assign intsink_metaReset = metaReset | intsink_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_33 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  RocketTile_metaAssert = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_33 <= 1'h0;
    end else if (reset) begin
      _T_33 <= 1'h0;
    end else begin
      _T_33 <= core_io_wfi;
    end
    if (metaReset) begin
      RocketTile_metaAssert <= 1'h0;
    end else begin
      RocketTile_metaAssert <= RocketTile_metaAssert | RocketTile_or0;
    end
  end
endmodule
module TLXbar_7(
  input         clock,
  input         reset,
  output        auto_in_1_a_ready,
  input         auto_in_1_a_valid,
  input  [31:0] auto_in_1_a_bits_address,
  output        auto_in_1_d_valid,
  output [2:0]  auto_in_1_d_bits_opcode,
  output [3:0]  auto_in_1_d_bits_size,
  output [63:0] auto_in_1_d_bits_data,
  output        auto_in_1_d_bits_corrupt,
  output        auto_in_0_a_ready,
  input         auto_in_0_a_valid,
  input  [2:0]  auto_in_0_a_bits_opcode,
  input  [2:0]  auto_in_0_a_bits_param,
  input  [3:0]  auto_in_0_a_bits_size,
  input         auto_in_0_a_bits_source,
  input  [31:0] auto_in_0_a_bits_address,
  input  [7:0]  auto_in_0_a_bits_mask,
  input  [63:0] auto_in_0_a_bits_data,
  input         auto_in_0_b_ready,
  output        auto_in_0_b_valid,
  output [1:0]  auto_in_0_b_bits_param,
  output [3:0]  auto_in_0_b_bits_size,
  output        auto_in_0_b_bits_source,
  output [31:0] auto_in_0_b_bits_address,
  output        auto_in_0_c_ready,
  input         auto_in_0_c_valid,
  input  [2:0]  auto_in_0_c_bits_opcode,
  input  [2:0]  auto_in_0_c_bits_param,
  input  [3:0]  auto_in_0_c_bits_size,
  input         auto_in_0_c_bits_source,
  input  [31:0] auto_in_0_c_bits_address,
  input  [63:0] auto_in_0_c_bits_data,
  input         auto_in_0_d_ready,
  output        auto_in_0_d_valid,
  output [2:0]  auto_in_0_d_bits_opcode,
  output [1:0]  auto_in_0_d_bits_param,
  output [3:0]  auto_in_0_d_bits_size,
  output        auto_in_0_d_bits_source,
  output [1:0]  auto_in_0_d_bits_sink,
  output        auto_in_0_d_bits_denied,
  output [63:0] auto_in_0_d_bits_data,
  output        auto_in_0_e_ready,
  input         auto_in_0_e_valid,
  input  [1:0]  auto_in_0_e_bits_sink,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [1:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_a_bits_corrupt,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [2:0]  auto_out_b_bits_opcode,
  input  [1:0]  auto_out_b_bits_param,
  input  [3:0]  auto_out_b_bits_size,
  input  [1:0]  auto_out_b_bits_source,
  input  [31:0] auto_out_b_bits_address,
  input  [7:0]  auto_out_b_bits_mask,
  input         auto_out_b_bits_corrupt,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [3:0]  auto_out_c_bits_size,
  output [1:0]  auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [3:0]  auto_out_d_bits_size,
  input  [1:0]  auto_out_d_bits_source,
  input  [1:0]  auto_out_d_bits_sink,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output [1:0]  auto_out_e_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         TLMonitor_halt,
  input         TLMonitor_1_halt
);
  wire  TLMonitor_clock; // @[Nodes.scala 25:25]
  wire  TLMonitor_reset; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_a_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_a_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_a_bits_opcode; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_a_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_a_bits_size; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_a_bits_source; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_io_in_a_bits_address; // @[Nodes.scala 25:25]
  wire [7:0] TLMonitor_io_in_a_bits_mask; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_b_bits_opcode; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_b_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_b_bits_size; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_bits_source; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_io_in_b_bits_address; // @[Nodes.scala 25:25]
  wire [7:0] TLMonitor_io_in_b_bits_mask; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_bits_corrupt; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_c_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_c_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_c_bits_opcode; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_c_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_c_bits_size; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_c_bits_source; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_io_in_c_bits_address; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_d_bits_opcode; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_d_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_d_bits_size; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_bits_source; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_d_bits_sink; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_bits_denied; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_bits_corrupt; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_e_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_e_valid; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_e_bits_sink; // @[Nodes.scala 25:25]
  wire [29:0] TLMonitor_io_covSum; // @[Nodes.scala 25:25]
  wire  TLMonitor_metaAssert; // @[Nodes.scala 25:25]
  wire  TLMonitor_metaReset; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_clock; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_reset; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_io_in_a_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_io_in_a_valid; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_1_io_in_a_bits_address; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_io_in_d_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_1_io_in_d_bits_opcode; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_1_io_in_d_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_1_io_in_d_bits_size; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_1_io_in_d_bits_sink; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_io_in_d_bits_denied; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_io_in_d_bits_corrupt; // @[Nodes.scala 25:25]
  wire [29:0] TLMonitor_1_io_covSum; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_metaAssert; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_metaReset; // @[Nodes.scala 25:25]
  wire  _T_59; // @[Parameters.scala 47:9]
  wire [26:0] _T_77; // @[package.scala 212:77]
  wire [8:0] _T_80; // @[Edges.scala 221:59]
  wire  _T_147; // @[Mux.scala 27:72]
  reg [8:0] _T_157; // @[Arbiter.scala 78:30]
  reg [31:0] _RAND_0;
  wire  _T_158; // @[Arbiter.scala 79:28]
  wire  _T_159; // @[Arbiter.scala 80:24]
  wire [1:0] _T_164; // @[Cat.scala 29:58]
  wire  _T_166; // @[Arbiter.scala 21:19]
  wire  _T_168; // @[Arbiter.scala 21:12]
  reg [1:0] _T_170; // @[Arbiter.scala 22:23]
  reg [31:0] _RAND_1;
  wire [1:0] _T_172; // @[Arbiter.scala 23:28]
  wire [3:0] _T_173; // @[Cat.scala 29:58]
  wire [3:0] _GEN_1; // @[package.scala 231:43]
  wire [3:0] _T_175; // @[package.scala 231:43]
  wire [3:0] _T_178; // @[Arbiter.scala 24:66]
  wire [3:0] _GEN_2; // @[Arbiter.scala 24:58]
  wire [3:0] _T_179; // @[Arbiter.scala 24:58]
  wire [1:0] _T_182; // @[Arbiter.scala 25:39]
  wire  _T_184; // @[Arbiter.scala 26:27]
  wire  _T_185; // @[Arbiter.scala 26:18]
  wire [1:0] _T_186; // @[Arbiter.scala 27:29]
  wire [2:0] _T_187; // @[package.scala 222:48]
  wire [1:0] _T_189; // @[package.scala 222:43]
  wire  _T_192; // @[Arbiter.scala 86:86]
  wire  _T_193; // @[Arbiter.scala 86:86]
  wire  _T_195; // @[Arbiter.scala 88:79]
  wire  _T_196; // @[Arbiter.scala 88:79]
  wire  _T_202; // @[Arbiter.scala 95:53]
  wire  _T_208; // @[Arbiter.scala 96:64]
  wire  _T_211; // @[Arbiter.scala 96:13]
  wire  _T_213; // @[Arbiter.scala 98:36]
  wire  _T_216; // @[Arbiter.scala 98:41]
  wire  _T_218; // @[Arbiter.scala 98:14]
  wire  _T_223; // @[Arbiter.scala 99:41]
  wire  _T_225; // @[Arbiter.scala 99:14]
  reg  _T_237_0; // @[Arbiter.scala 107:26]
  reg [31:0] _RAND_2;
  wire  _T_238_0; // @[Arbiter.scala 108:30]
  reg  _T_237_1; // @[Arbiter.scala 107:26]
  reg [31:0] _RAND_3;
  wire  _T_238_1; // @[Arbiter.scala 108:30]
  wire  _T_244; // @[Mux.scala 27:72]
  wire  _T_245; // @[Mux.scala 27:72]
  wire  _T_246; // @[Mux.scala 27:72]
  wire  _T_248; // @[Arbiter.scala 116:29]
  wire  _T_232; // @[ReadyValidCancel.scala 52:33]
  wire [8:0] _GEN_3; // @[Arbiter.scala 104:52]
  wire [8:0] _T_234; // @[Arbiter.scala 104:52]
  wire  _T_240_0; // @[Arbiter.scala 112:24]
  wire  _T_240_1; // @[Arbiter.scala 112:24]
  wire [1:0] _T_9_0_a_bits_source; // @[Xbar.scala 225:18 BundleMap.scala 248:19 Xbar.scala 231:29]
  wire [116:0] _T_259; // @[Mux.scala 27:72]
  wire [116:0] _T_260; // @[Mux.scala 27:72]
  wire [116:0] _T_267; // @[Mux.scala 27:72]
  wire [116:0] _T_268; // @[Mux.scala 27:72]
  wire [116:0] _T_269; // @[Mux.scala 27:72]
  reg [2:0] TLXbar_7_state; // @[Register tracking TLXbar_7 state]
  reg [31:0] _RAND_4;
  reg  TLXbar_7_cov [0:7]; // @[Coverage map for TLXbar_7]
  reg [31:0] _RAND_5;
  wire  TLXbar_7_cov_read_data; // @[Coverage map for TLXbar_7]
  wire [2:0] TLXbar_7_cov_read_addr; // @[Coverage map for TLXbar_7]
  wire  TLXbar_7_cov_write_data; // @[Coverage map for TLXbar_7]
  wire [2:0] TLXbar_7_cov_write_addr; // @[Coverage map for TLXbar_7]
  wire  TLXbar_7_cov_write_mask; // @[Coverage map for TLXbar_7]
  wire  TLXbar_7_cov_write_en; // @[Coverage map for TLXbar_7]
  reg [29:0] TLXbar_7_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_6;
  wire [1:0] _T_170_shl;
  wire [2:0] _T_170_pad;
  wire [2:0] _T_237_0_shl;
  wire [2:0] _T_237_0_pad;
  wire [2:0] _T_237_1_shl;
  wire [2:0] _T_237_1_pad;
  wire [2:0] TLXbar_7_xor2;
  wire [2:0] TLXbar_7_xor0;
  wire [29:0] TLMonitor_sum;
  wire [29:0] TLMonitor_1_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  TLMonitor_metaAssert_wire;
  wire  TLMonitor_1_metaAssert_wire;
  wire  TLXbar_7_or4;
  wire  TLXbar_7_or1;
  wire  TLXbar_7_or6;
  wire  TLXbar_7_or2;
  wire  TLXbar_7_or0;
  reg  TLXbar_7_metaAssert;
  reg [31:0] _RAND_7;
  TLMonitor_35 TLMonitor ( // @[Nodes.scala 25:25]
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_b_ready(TLMonitor_io_in_b_ready),
    .io_in_b_valid(TLMonitor_io_in_b_valid),
    .io_in_b_bits_opcode(TLMonitor_io_in_b_bits_opcode),
    .io_in_b_bits_param(TLMonitor_io_in_b_bits_param),
    .io_in_b_bits_size(TLMonitor_io_in_b_bits_size),
    .io_in_b_bits_source(TLMonitor_io_in_b_bits_source),
    .io_in_b_bits_address(TLMonitor_io_in_b_bits_address),
    .io_in_b_bits_mask(TLMonitor_io_in_b_bits_mask),
    .io_in_b_bits_corrupt(TLMonitor_io_in_b_bits_corrupt),
    .io_in_c_ready(TLMonitor_io_in_c_ready),
    .io_in_c_valid(TLMonitor_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_io_in_c_bits_address),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt),
    .io_in_e_ready(TLMonitor_io_in_e_ready),
    .io_in_e_valid(TLMonitor_io_in_e_valid),
    .io_in_e_bits_sink(TLMonitor_io_in_e_bits_sink),
    .io_covSum(TLMonitor_io_covSum),
    .metaAssert(TLMonitor_metaAssert),
    .metaReset(TLMonitor_metaReset)
  );
  TLMonitor_36 TLMonitor_1 ( // @[Nodes.scala 25:25]
    .clock(TLMonitor_1_clock),
    .reset(TLMonitor_1_reset),
    .io_in_a_ready(TLMonitor_1_io_in_a_ready),
    .io_in_a_valid(TLMonitor_1_io_in_a_valid),
    .io_in_a_bits_address(TLMonitor_1_io_in_a_bits_address),
    .io_in_d_valid(TLMonitor_1_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_1_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_1_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_1_io_in_d_bits_size),
    .io_in_d_bits_sink(TLMonitor_1_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_1_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_1_io_in_d_bits_corrupt),
    .io_covSum(TLMonitor_1_io_covSum),
    .metaAssert(TLMonitor_1_metaAssert),
    .metaReset(TLMonitor_1_metaReset)
  );
  assign _T_59 = auto_out_d_bits_source == 2'h2; // @[Parameters.scala 47:9]
  assign _T_77 = 27'hfff << auto_in_0_a_bits_size; // @[package.scala 212:77]
  assign _T_80 = ~_T_77[11:3]; // @[Edges.scala 221:59]
  assign _T_147 = ~auto_out_d_bits_source[1] & auto_in_0_d_ready; // @[Mux.scala 27:72]
  assign _T_158 = _T_157 == 9'h0; // @[Arbiter.scala 79:28]
  assign _T_159 = _T_158 & auto_out_a_ready; // @[Arbiter.scala 80:24]
  assign _T_164 = {auto_in_1_a_valid,auto_in_0_a_valid}; // @[Cat.scala 29:58]
  assign _T_166 = _T_164 == _T_164; // @[Arbiter.scala 21:19]
  assign _T_168 = _T_166 | reset; // @[Arbiter.scala 21:12]
  assign _T_172 = _T_164 & ~_T_170; // @[Arbiter.scala 23:28]
  assign _T_173 = {_T_172,auto_in_1_a_valid,auto_in_0_a_valid}; // @[Cat.scala 29:58]
  assign _GEN_1 = {{1'd0}, _T_173[3:1]}; // @[package.scala 231:43]
  assign _T_175 = _T_173 | _GEN_1; // @[package.scala 231:43]
  assign _T_178 = {_T_170, 2'h0}; // @[Arbiter.scala 24:66]
  assign _GEN_2 = {{1'd0}, _T_175[3:1]}; // @[Arbiter.scala 24:58]
  assign _T_179 = _GEN_2 | _T_178; // @[Arbiter.scala 24:58]
  assign _T_182 = _T_179[3:2] & _T_179[1:0]; // @[Arbiter.scala 25:39]
  assign _T_184 = |_T_164; // @[Arbiter.scala 26:27]
  assign _T_185 = _T_159 & _T_184; // @[Arbiter.scala 26:18]
  assign _T_186 = ~_T_182 & _T_164; // @[Arbiter.scala 27:29]
  assign _T_187 = {_T_186, 1'h0}; // @[package.scala 222:48]
  assign _T_189 = _T_186 | _T_187[1:0]; // @[package.scala 222:43]
  assign _T_192 = ~_T_182[0]; // @[Arbiter.scala 86:86]
  assign _T_193 = ~_T_182[1]; // @[Arbiter.scala 86:86]
  assign _T_195 = _T_192 & auto_in_0_a_valid; // @[Arbiter.scala 88:79]
  assign _T_196 = _T_193 & auto_in_1_a_valid; // @[Arbiter.scala 88:79]
  assign _T_202 = _T_195 | _T_196; // @[Arbiter.scala 95:53]
  assign _T_208 = ~_T_195 | ~_T_196; // @[Arbiter.scala 96:64]
  assign _T_211 = _T_208 | reset; // @[Arbiter.scala 96:13]
  assign _T_213 = auto_in_0_a_valid | auto_in_1_a_valid; // @[Arbiter.scala 98:36]
  assign _T_216 = ~_T_213 | _T_202; // @[Arbiter.scala 98:41]
  assign _T_218 = _T_216 | reset; // @[Arbiter.scala 98:14]
  assign _T_223 = ~_T_213 | _T_213; // @[Arbiter.scala 99:41]
  assign _T_225 = _T_223 | reset; // @[Arbiter.scala 99:14]
  assign _T_238_0 = _T_158 ? _T_195 : _T_237_0; // @[Arbiter.scala 108:30]
  assign _T_238_1 = _T_158 ? _T_196 : _T_237_1; // @[Arbiter.scala 108:30]
  assign _T_244 = _T_237_0 & auto_in_0_a_valid; // @[Mux.scala 27:72]
  assign _T_245 = _T_237_1 & auto_in_1_a_valid; // @[Mux.scala 27:72]
  assign _T_246 = _T_244 | _T_245; // @[Mux.scala 27:72]
  assign _T_248 = _T_158 ? _T_213 : _T_246; // @[Arbiter.scala 116:29]
  assign _T_232 = auto_out_a_ready & _T_248; // @[ReadyValidCancel.scala 52:33]
  assign _GEN_3 = {{8'd0}, _T_232}; // @[Arbiter.scala 104:52]
  assign _T_234 = _T_157 - _GEN_3; // @[Arbiter.scala 104:52]
  assign _T_240_0 = _T_158 ? _T_192 : _T_237_0; // @[Arbiter.scala 112:24]
  assign _T_240_1 = _T_158 ? _T_193 : _T_237_1; // @[Arbiter.scala 112:24]
  assign _T_9_0_a_bits_source = {{1'd0}, auto_in_0_a_bits_source}; // @[Xbar.scala 225:18 BundleMap.scala 248:19 Xbar.scala 231:29]
  assign _T_259 = {auto_in_0_a_bits_opcode,auto_in_0_a_bits_param,auto_in_0_a_bits_size,_T_9_0_a_bits_source,auto_in_0_a_bits_address,auto_in_0_a_bits_mask,auto_in_0_a_bits_data,1'h0}; // @[Mux.scala 27:72]
  assign _T_260 = _T_238_0 ? _T_259 : 117'h0; // @[Mux.scala 27:72]
  assign _T_267 = {12'h81a,auto_in_1_a_bits_address,8'hff,65'h0}; // @[Mux.scala 27:72]
  assign _T_268 = _T_238_1 ? _T_267 : 117'h0; // @[Mux.scala 27:72]
  assign _T_269 = _T_260 | _T_268; // @[Mux.scala 27:72]
  assign auto_in_1_a_ready = auto_out_a_ready & _T_240_1; // @[LazyModule.scala 303:16]
  assign auto_in_1_d_valid = auto_out_d_valid & _T_59; // @[LazyModule.scala 303:16]
  assign auto_in_1_d_bits_opcode = auto_out_d_bits_opcode; // @[LazyModule.scala 303:16]
  assign auto_in_1_d_bits_size = auto_out_d_bits_size; // @[LazyModule.scala 303:16]
  assign auto_in_1_d_bits_data = auto_out_d_bits_data; // @[LazyModule.scala 303:16]
  assign auto_in_1_d_bits_corrupt = auto_out_d_bits_corrupt; // @[LazyModule.scala 303:16]
  assign auto_in_0_a_ready = auto_out_a_ready & _T_240_0; // @[LazyModule.scala 303:16]
  assign auto_in_0_b_valid = auto_out_b_valid & ~auto_out_b_bits_source[1]; // @[LazyModule.scala 303:16]
  assign auto_in_0_b_bits_param = auto_out_b_bits_param; // @[LazyModule.scala 303:16]
  assign auto_in_0_b_bits_size = auto_out_b_bits_size; // @[LazyModule.scala 303:16]
  assign auto_in_0_b_bits_source = auto_out_b_bits_source[0]; // @[LazyModule.scala 303:16]
  assign auto_in_0_b_bits_address = auto_out_b_bits_address; // @[LazyModule.scala 303:16]
  assign auto_in_0_c_ready = auto_out_c_ready; // @[LazyModule.scala 303:16]
  assign auto_in_0_d_valid = auto_out_d_valid & ~auto_out_d_bits_source[1]; // @[LazyModule.scala 303:16]
  assign auto_in_0_d_bits_opcode = auto_out_d_bits_opcode; // @[LazyModule.scala 303:16]
  assign auto_in_0_d_bits_param = auto_out_d_bits_param; // @[LazyModule.scala 303:16]
  assign auto_in_0_d_bits_size = auto_out_d_bits_size; // @[LazyModule.scala 303:16]
  assign auto_in_0_d_bits_source = auto_out_d_bits_source[0]; // @[LazyModule.scala 303:16]
  assign auto_in_0_d_bits_sink = auto_out_d_bits_sink; // @[LazyModule.scala 303:16]
  assign auto_in_0_d_bits_denied = auto_out_d_bits_denied; // @[LazyModule.scala 303:16]
  assign auto_in_0_d_bits_data = auto_out_d_bits_data; // @[LazyModule.scala 303:16]
  assign auto_in_0_e_ready = auto_out_e_ready; // @[LazyModule.scala 303:16]
  assign auto_out_a_valid = _T_158 ? _T_213 : _T_246; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_opcode = _T_269[116:114]; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_param = _T_269[113:111]; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_size = _T_269[110:107]; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_source = _T_269[106:105]; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_address = _T_269[104:73]; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_mask = _T_269[72:65]; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_data = _T_269[64:1]; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_corrupt = _T_269[0]; // @[LazyModule.scala 305:12]
  assign auto_out_b_ready = ~auto_out_b_bits_source[1] & auto_in_0_b_ready; // @[LazyModule.scala 305:12]
  assign auto_out_c_valid = auto_in_0_c_valid; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_opcode = auto_in_0_c_bits_opcode; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_param = auto_in_0_c_bits_param; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_size = auto_in_0_c_bits_size; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_source = {{1'd0}, auto_in_0_c_bits_source}; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_address = auto_in_0_c_bits_address; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_data = auto_in_0_c_bits_data; // @[LazyModule.scala 305:12]
  assign auto_out_d_ready = _T_147 | _T_59; // @[LazyModule.scala 305:12]
  assign auto_out_e_valid = auto_in_0_e_valid; // @[LazyModule.scala 305:12]
  assign auto_out_e_bits_sink = auto_in_0_e_bits_sink; // @[LazyModule.scala 305:12]
  assign TLMonitor_clock = clock;
  assign TLMonitor_reset = reset;
  assign TLMonitor_io_in_a_ready = auto_out_a_ready & _T_240_0; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_valid = auto_in_0_a_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_opcode = auto_in_0_a_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_param = auto_in_0_a_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_size = auto_in_0_a_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_source = auto_in_0_a_bits_source; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_address = auto_in_0_a_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_mask = auto_in_0_a_bits_mask; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_ready = auto_in_0_b_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_valid = auto_out_b_valid & ~auto_out_b_bits_source[1]; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_opcode = auto_out_b_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_param = auto_out_b_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_size = auto_out_b_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_source = auto_out_b_bits_source[0]; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_address = auto_out_b_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_mask = auto_out_b_bits_mask; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_corrupt = auto_out_b_bits_corrupt; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_ready = auto_out_c_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_valid = auto_in_0_c_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_opcode = auto_in_0_c_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_param = auto_in_0_c_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_size = auto_in_0_c_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_source = auto_in_0_c_bits_source; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_address = auto_in_0_c_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_ready = auto_in_0_d_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_valid = auto_out_d_valid & ~auto_out_d_bits_source[1]; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_source = auto_out_d_bits_source[0]; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_e_ready = auto_out_e_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_e_valid = auto_in_0_e_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_e_bits_sink = auto_in_0_e_bits_sink; // @[Nodes.scala 26:19]
  assign TLMonitor_1_clock = clock;
  assign TLMonitor_1_reset = reset;
  assign TLMonitor_1_io_in_a_ready = auto_out_a_ready & _T_240_1; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_a_valid = auto_in_1_a_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_a_bits_address = auto_in_1_a_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_valid = auto_out_d_valid & _T_59; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 26:19]
  assign TLXbar_7_cov_read_addr = TLXbar_7_state;
  assign TLXbar_7_cov_read_data = TLXbar_7_cov[TLXbar_7_cov_read_addr]; // @[Coverage map for TLXbar_7]
  assign TLXbar_7_cov_write_data = 1'h1;
  assign TLXbar_7_cov_write_addr = TLXbar_7_state;
  assign TLXbar_7_cov_write_mask = 1'h1;
  assign TLXbar_7_cov_write_en = 1'h1;
  assign _T_170_shl = _T_170;
  assign _T_170_pad = {1'h0,_T_170_shl};
  assign _T_237_0_shl = {_T_237_0, 2'h0};
  assign _T_237_0_pad = _T_237_0_shl;
  assign _T_237_1_shl = {_T_237_1, 2'h0};
  assign _T_237_1_pad = _T_237_1_shl;
  assign TLXbar_7_xor2 = _T_237_0_pad ^ _T_237_1_pad;
  assign TLXbar_7_xor0 = _T_170_pad ^ TLXbar_7_xor2;
  assign TLMonitor_sum = TLXbar_7_covSum + TLMonitor_io_covSum;
  assign TLMonitor_1_sum = TLMonitor_sum + TLMonitor_1_io_covSum;
  assign io_covSum = TLMonitor_1_sum;
  assign stopEn0 = ~_T_168;
  assign stopEn1 = ~_T_211;
  assign stopEn2 = ~_T_218;
  assign stopEn3 = ~_T_225;
  assign TLMonitor_metaAssert_wire = TLMonitor_metaAssert;
  assign TLMonitor_1_metaAssert_wire = TLMonitor_1_metaAssert;
  assign TLXbar_7_or4 = stopEn1 | stopEn2;
  assign TLXbar_7_or1 = stopEn0 | TLXbar_7_or4;
  assign TLXbar_7_or6 = TLMonitor_metaAssert_wire | TLMonitor_1_metaAssert_wire;
  assign TLXbar_7_or2 = stopEn3 | TLXbar_7_or6;
  assign TLXbar_7_or0 = TLXbar_7_or1 | TLXbar_7_or2;
  assign metaAssert = TLXbar_7_metaAssert;
  assign TLMonitor_metaReset = metaReset | TLMonitor_halt;
  assign TLMonitor_1_metaReset = metaReset | TLMonitor_1_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_157 = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_170 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_237_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_237_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  TLXbar_7_state = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    TLXbar_7_cov[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  TLXbar_7_covSum = _RAND_6[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  TLXbar_7_metaAssert = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_157 <= 9'h0;
    end else if (reset) begin
      _T_157 <= 9'h0;
    end else if (_T_159) begin
      if (_T_195) begin
        if (~auto_in_0_a_bits_opcode[2]) begin
          _T_157 <= _T_80;
        end else begin
          _T_157 <= 9'h0;
        end
      end else begin
        _T_157 <= 9'h0;
      end
    end else begin
      _T_157 <= _T_234;
    end
    if (metaReset) begin
      _T_170 <= 2'h0;
    end else if (reset) begin
      _T_170 <= 2'h3;
    end else if (_T_185) begin
      _T_170 <= _T_189;
    end
    if (metaReset) begin
      _T_237_0 <= 1'h0;
    end else if (reset) begin
      _T_237_0 <= 1'h0;
    end else if (_T_158) begin
      _T_237_0 <= _T_195;
    end
    if (metaReset) begin
      _T_237_1 <= 1'h0;
    end else if (reset) begin
      _T_237_1 <= 1'h0;
    end else if (_T_158) begin
      _T_237_1 <= _T_196;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_168) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:21 assert (valid === valids)\n"); // @[Arbiter.scala 21:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_168) begin
          $fatal; // @[Arbiter.scala 21:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_211) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:96 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Arbiter.scala 96:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_211) begin
          $fatal; // @[Arbiter.scala 96:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_218) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:98 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"); // @[Arbiter.scala 98:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_218) begin
          $fatal; // @[Arbiter.scala 98:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_225) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:99 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"); // @[Arbiter.scala 99:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_225) begin
          $fatal; // @[Arbiter.scala 99:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    TLXbar_7_state <= TLXbar_7_xor0;
    if (!(TLXbar_7_cov_read_data)) begin
      TLXbar_7_covSum <= TLXbar_7_covSum + 1'h1;
    end
    if (metaReset) begin
      TLXbar_7_metaAssert <= 1'h0;
    end else begin
      TLXbar_7_metaAssert <= TLXbar_7_metaAssert | TLXbar_7_or0;
    end
  end
  always @(posedge clock) begin
    if(TLXbar_7_cov_write_en & TLXbar_7_cov_write_mask) begin
      TLXbar_7_cov[TLXbar_7_cov_write_addr] <= TLXbar_7_cov_write_data; // @[Coverage map for TLXbar_7]
    end
  end
endmodule
module IntXbar_1(
  input         auto_int_in_3_0,
  input         auto_int_in_2_0,
  input         auto_int_in_1_0,
  input         auto_int_in_1_1,
  input         auto_int_in_0_0,
  output        auto_int_out_0,
  output        auto_int_out_1,
  output        auto_int_out_2,
  output        auto_int_out_3,
  output        auto_int_out_4,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] IntXbar_1_covSum;
  assign auto_int_out_0 = auto_int_in_0_0; // @[LazyModule.scala 305:12]
  assign auto_int_out_1 = auto_int_in_1_0; // @[LazyModule.scala 305:12]
  assign auto_int_out_2 = auto_int_in_1_1; // @[LazyModule.scala 305:12]
  assign auto_int_out_3 = auto_int_in_2_0; // @[LazyModule.scala 305:12]
  assign auto_int_out_4 = auto_int_in_3_0; // @[LazyModule.scala 305:12]
  assign IntXbar_1_covSum = 30'h0;
  assign io_covSum = IntXbar_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module BundleBridgeNexus(
  input         auto_in,
  output        auto_out_0,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] BundleBridgeNexus_covSum;
  assign auto_out_0 = auto_in; // @[LazyModule.scala 305:12]
  assign BundleBridgeNexus_covSum = 30'h0;
  assign io_covSum = BundleBridgeNexus_covSum;
  assign metaAssert = 1'h0;
endmodule
module BundleBridgeNexus_1(
  input  [31:0] auto_in,
  output [31:0] auto_out_1,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] BundleBridgeNexus_1_covSum;
  assign auto_out_1 = auto_in; // @[LazyModule.scala 305:12]
  assign BundleBridgeNexus_1_covSum = 30'h0;
  assign io_covSum = BundleBridgeNexus_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module DCache(
  input         gated_clock,
  input         reset,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output        auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [1:0]  auto_out_b_bits_param,
  input  [3:0]  auto_out_b_bits_size,
  input         auto_out_b_bits_source,
  input  [31:0] auto_out_b_bits_address,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [3:0]  auto_out_c_bits_size,
  output        auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [3:0]  auto_out_d_bits_size,
  input         auto_out_d_bits_source,
  input  [1:0]  auto_out_d_bits_sink,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output [1:0]  auto_out_e_bits_sink,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_addr,
  input  [6:0]  io_cpu_req_bits_tag,
  input  [4:0]  io_cpu_req_bits_cmd,
  input  [1:0]  io_cpu_req_bits_size,
  input         io_cpu_req_bits_signed,
  input         io_cpu_req_bits_phys,
  input         io_cpu_s1_kill,
  input  [63:0] io_cpu_s1_data_data,
  output        io_cpu_s2_nack,
  output        io_cpu_resp_valid,
  output [6:0]  io_cpu_resp_bits_tag,
  output [1:0]  io_cpu_resp_bits_size,
  output [63:0] io_cpu_resp_bits_data,
  output        io_cpu_resp_bits_replay,
  output        io_cpu_resp_bits_has_data,
  output [63:0] io_cpu_resp_bits_data_word_bypass,
  output        io_cpu_replay_next,
  output        io_cpu_s2_xcpt_ma_ld,
  output        io_cpu_s2_xcpt_ma_st,
  output        io_cpu_s2_xcpt_pf_ld,
  output        io_cpu_s2_xcpt_pf_st,
  output        io_cpu_s2_xcpt_ae_ld,
  output        io_cpu_s2_xcpt_ae_st,
  output        io_cpu_ordered,
  output        io_cpu_perf_release,
  output        io_cpu_perf_grant,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input         io_ptw_status_debug,
  input  [1:0]  io_ptw_status_dprv,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         MaxPeriodFibonacciLFSR_halt,
  input         pma_checker_halt,
  input         tlb_halt,
  input         data_halt,
  output [19:0] Checking_DCache_regstate,	//Jaewon_DCache_regstate
  output [29:0] Checking_DCache_covSum	//Jaewon_DCache_regstate
  );
  assign Checking_DCache_regstate = DCache_state; 	//Jaewon_DCache_regstate
  assign Checking_DCache_covSum = DCache_covSum; 	//Jaewon_DCache_regstate
  wire  tlb_clock; // @[DCache.scala 115:19]
  wire  tlb_reset; // @[DCache.scala 115:19]
  wire  tlb_io_req_ready; // @[DCache.scala 115:19]
  wire  tlb_io_req_valid; // @[DCache.scala 115:19]
  wire [39:0] tlb_io_req_bits_vaddr; // @[DCache.scala 115:19]
  wire  tlb_io_req_bits_passthrough; // @[DCache.scala 115:19]
  wire [1:0] tlb_io_req_bits_size; // @[DCache.scala 115:19]
  wire [4:0] tlb_io_req_bits_cmd; // @[DCache.scala 115:19]
  wire  tlb_io_resp_miss; // @[DCache.scala 115:19]
  wire [31:0] tlb_io_resp_paddr; // @[DCache.scala 115:19]
  wire  tlb_io_resp_pf_ld; // @[DCache.scala 115:19]
  wire  tlb_io_resp_pf_st; // @[DCache.scala 115:19]
  wire  tlb_io_resp_ae_ld; // @[DCache.scala 115:19]
  wire  tlb_io_resp_ae_st; // @[DCache.scala 115:19]
  wire  tlb_io_resp_ma_ld; // @[DCache.scala 115:19]
  wire  tlb_io_resp_ma_st; // @[DCache.scala 115:19]
  wire  tlb_io_resp_cacheable; // @[DCache.scala 115:19]
  wire  tlb_io_sfence_valid; // @[DCache.scala 115:19]
  wire  tlb_io_sfence_bits_rs1; // @[DCache.scala 115:19]
  wire  tlb_io_sfence_bits_rs2; // @[DCache.scala 115:19]
  wire [38:0] tlb_io_sfence_bits_addr; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_req_ready; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_req_valid; // @[DCache.scala 115:19]
  wire [26:0] tlb_io_ptw_req_bits_bits_addr; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_resp_valid; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_resp_bits_ae; // @[DCache.scala 115:19]
  wire [53:0] tlb_io_ptw_resp_bits_pte_ppn; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_resp_bits_pte_d; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_resp_bits_pte_a; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_resp_bits_pte_g; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_resp_bits_pte_u; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_resp_bits_pte_x; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_resp_bits_pte_w; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_resp_bits_pte_r; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_resp_bits_pte_v; // @[DCache.scala 115:19]
  wire [1:0] tlb_io_ptw_resp_bits_level; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_resp_bits_homogeneous; // @[DCache.scala 115:19]
  wire [3:0] tlb_io_ptw_ptbr_mode; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_status_debug; // @[DCache.scala 115:19]
  wire [1:0] tlb_io_ptw_status_dprv; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_status_mxr; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_status_sum; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_0_cfg_l; // @[DCache.scala 115:19]
  wire [1:0] tlb_io_ptw_pmp_0_cfg_a; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_0_cfg_x; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_0_cfg_w; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_0_cfg_r; // @[DCache.scala 115:19]
  wire [29:0] tlb_io_ptw_pmp_0_addr; // @[DCache.scala 115:19]
  wire [31:0] tlb_io_ptw_pmp_0_mask; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_1_cfg_l; // @[DCache.scala 115:19]
  wire [1:0] tlb_io_ptw_pmp_1_cfg_a; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_1_cfg_x; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_1_cfg_w; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_1_cfg_r; // @[DCache.scala 115:19]
  wire [29:0] tlb_io_ptw_pmp_1_addr; // @[DCache.scala 115:19]
  wire [31:0] tlb_io_ptw_pmp_1_mask; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_2_cfg_l; // @[DCache.scala 115:19]
  wire [1:0] tlb_io_ptw_pmp_2_cfg_a; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_2_cfg_x; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_2_cfg_w; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_2_cfg_r; // @[DCache.scala 115:19]
  wire [29:0] tlb_io_ptw_pmp_2_addr; // @[DCache.scala 115:19]
  wire [31:0] tlb_io_ptw_pmp_2_mask; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_3_cfg_l; // @[DCache.scala 115:19]
  wire [1:0] tlb_io_ptw_pmp_3_cfg_a; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_3_cfg_x; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_3_cfg_w; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_3_cfg_r; // @[DCache.scala 115:19]
  wire [29:0] tlb_io_ptw_pmp_3_addr; // @[DCache.scala 115:19]
  wire [31:0] tlb_io_ptw_pmp_3_mask; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_4_cfg_l; // @[DCache.scala 115:19]
  wire [1:0] tlb_io_ptw_pmp_4_cfg_a; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_4_cfg_x; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_4_cfg_w; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_4_cfg_r; // @[DCache.scala 115:19]
  wire [29:0] tlb_io_ptw_pmp_4_addr; // @[DCache.scala 115:19]
  wire [31:0] tlb_io_ptw_pmp_4_mask; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_5_cfg_l; // @[DCache.scala 115:19]
  wire [1:0] tlb_io_ptw_pmp_5_cfg_a; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_5_cfg_x; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_5_cfg_w; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_5_cfg_r; // @[DCache.scala 115:19]
  wire [29:0] tlb_io_ptw_pmp_5_addr; // @[DCache.scala 115:19]
  wire [31:0] tlb_io_ptw_pmp_5_mask; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_6_cfg_l; // @[DCache.scala 115:19]
  wire [1:0] tlb_io_ptw_pmp_6_cfg_a; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_6_cfg_x; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_6_cfg_w; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_6_cfg_r; // @[DCache.scala 115:19]
  wire [29:0] tlb_io_ptw_pmp_6_addr; // @[DCache.scala 115:19]
  wire [31:0] tlb_io_ptw_pmp_6_mask; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_7_cfg_l; // @[DCache.scala 115:19]
  wire [1:0] tlb_io_ptw_pmp_7_cfg_a; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_7_cfg_x; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_7_cfg_w; // @[DCache.scala 115:19]
  wire  tlb_io_ptw_pmp_7_cfg_r; // @[DCache.scala 115:19]
  wire [29:0] tlb_io_ptw_pmp_7_addr; // @[DCache.scala 115:19]
  wire [31:0] tlb_io_ptw_pmp_7_mask; // @[DCache.scala 115:19]
  wire [29:0] tlb_io_covSum; // @[DCache.scala 115:19]
  wire  tlb_metaAssert; // @[DCache.scala 115:19]
  wire  tlb_metaReset; // @[DCache.scala 115:19]
  wire  pma_checker_clock; // @[DCache.scala 116:27]
  wire  pma_checker_reset; // @[DCache.scala 116:27]
  wire  pma_checker_io_req_ready; // @[DCache.scala 116:27]
  wire  pma_checker_io_req_valid; // @[DCache.scala 116:27]
  wire [39:0] pma_checker_io_req_bits_vaddr; // @[DCache.scala 116:27]
  wire  pma_checker_io_req_bits_passthrough; // @[DCache.scala 116:27]
  wire [1:0] pma_checker_io_req_bits_size; // @[DCache.scala 116:27]
  wire [4:0] pma_checker_io_req_bits_cmd; // @[DCache.scala 116:27]
  wire  pma_checker_io_resp_miss; // @[DCache.scala 116:27]
  wire [31:0] pma_checker_io_resp_paddr; // @[DCache.scala 116:27]
  wire  pma_checker_io_resp_pf_ld; // @[DCache.scala 116:27]
  wire  pma_checker_io_resp_pf_st; // @[DCache.scala 116:27]
  wire  pma_checker_io_resp_ae_ld; // @[DCache.scala 116:27]
  wire  pma_checker_io_resp_ae_st; // @[DCache.scala 116:27]
  wire  pma_checker_io_resp_ma_ld; // @[DCache.scala 116:27]
  wire  pma_checker_io_resp_ma_st; // @[DCache.scala 116:27]
  wire  pma_checker_io_resp_cacheable; // @[DCache.scala 116:27]
  wire  pma_checker_io_sfence_valid; // @[DCache.scala 116:27]
  wire  pma_checker_io_sfence_bits_rs1; // @[DCache.scala 116:27]
  wire  pma_checker_io_sfence_bits_rs2; // @[DCache.scala 116:27]
  wire [38:0] pma_checker_io_sfence_bits_addr; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_req_ready; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_req_valid; // @[DCache.scala 116:27]
  wire [26:0] pma_checker_io_ptw_req_bits_bits_addr; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_resp_valid; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_resp_bits_ae; // @[DCache.scala 116:27]
  wire [53:0] pma_checker_io_ptw_resp_bits_pte_ppn; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_resp_bits_pte_d; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_resp_bits_pte_a; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_resp_bits_pte_g; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_resp_bits_pte_u; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_resp_bits_pte_x; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_resp_bits_pte_w; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_resp_bits_pte_r; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_resp_bits_pte_v; // @[DCache.scala 116:27]
  wire [1:0] pma_checker_io_ptw_resp_bits_level; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_resp_bits_homogeneous; // @[DCache.scala 116:27]
  wire [3:0] pma_checker_io_ptw_ptbr_mode; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_status_debug; // @[DCache.scala 116:27]
  wire [1:0] pma_checker_io_ptw_status_dprv; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_status_mxr; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_status_sum; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_0_cfg_l; // @[DCache.scala 116:27]
  wire [1:0] pma_checker_io_ptw_pmp_0_cfg_a; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_0_cfg_x; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_0_cfg_w; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_0_cfg_r; // @[DCache.scala 116:27]
  wire [29:0] pma_checker_io_ptw_pmp_0_addr; // @[DCache.scala 116:27]
  wire [31:0] pma_checker_io_ptw_pmp_0_mask; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_1_cfg_l; // @[DCache.scala 116:27]
  wire [1:0] pma_checker_io_ptw_pmp_1_cfg_a; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_1_cfg_x; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_1_cfg_w; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_1_cfg_r; // @[DCache.scala 116:27]
  wire [29:0] pma_checker_io_ptw_pmp_1_addr; // @[DCache.scala 116:27]
  wire [31:0] pma_checker_io_ptw_pmp_1_mask; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_2_cfg_l; // @[DCache.scala 116:27]
  wire [1:0] pma_checker_io_ptw_pmp_2_cfg_a; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_2_cfg_x; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_2_cfg_w; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_2_cfg_r; // @[DCache.scala 116:27]
  wire [29:0] pma_checker_io_ptw_pmp_2_addr; // @[DCache.scala 116:27]
  wire [31:0] pma_checker_io_ptw_pmp_2_mask; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_3_cfg_l; // @[DCache.scala 116:27]
  wire [1:0] pma_checker_io_ptw_pmp_3_cfg_a; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_3_cfg_x; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_3_cfg_w; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_3_cfg_r; // @[DCache.scala 116:27]
  wire [29:0] pma_checker_io_ptw_pmp_3_addr; // @[DCache.scala 116:27]
  wire [31:0] pma_checker_io_ptw_pmp_3_mask; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_4_cfg_l; // @[DCache.scala 116:27]
  wire [1:0] pma_checker_io_ptw_pmp_4_cfg_a; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_4_cfg_x; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_4_cfg_w; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_4_cfg_r; // @[DCache.scala 116:27]
  wire [29:0] pma_checker_io_ptw_pmp_4_addr; // @[DCache.scala 116:27]
  wire [31:0] pma_checker_io_ptw_pmp_4_mask; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_5_cfg_l; // @[DCache.scala 116:27]
  wire [1:0] pma_checker_io_ptw_pmp_5_cfg_a; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_5_cfg_x; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_5_cfg_w; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_5_cfg_r; // @[DCache.scala 116:27]
  wire [29:0] pma_checker_io_ptw_pmp_5_addr; // @[DCache.scala 116:27]
  wire [31:0] pma_checker_io_ptw_pmp_5_mask; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_6_cfg_l; // @[DCache.scala 116:27]
  wire [1:0] pma_checker_io_ptw_pmp_6_cfg_a; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_6_cfg_x; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_6_cfg_w; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_6_cfg_r; // @[DCache.scala 116:27]
  wire [29:0] pma_checker_io_ptw_pmp_6_addr; // @[DCache.scala 116:27]
  wire [31:0] pma_checker_io_ptw_pmp_6_mask; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_7_cfg_l; // @[DCache.scala 116:27]
  wire [1:0] pma_checker_io_ptw_pmp_7_cfg_a; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_7_cfg_x; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_7_cfg_w; // @[DCache.scala 116:27]
  wire  pma_checker_io_ptw_pmp_7_cfg_r; // @[DCache.scala 116:27]
  wire [29:0] pma_checker_io_ptw_pmp_7_addr; // @[DCache.scala 116:27]
  wire [31:0] pma_checker_io_ptw_pmp_7_mask; // @[DCache.scala 116:27]
  wire [29:0] pma_checker_io_covSum; // @[DCache.scala 116:27]
  wire  pma_checker_metaAssert; // @[DCache.scala 116:27]
  wire  pma_checker_metaReset; // @[DCache.scala 116:27]
  wire  MaxPeriodFibonacciLFSR_clock; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_reset; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_increment; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_0; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_1; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_2; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_3; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_4; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_5; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_6; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_7; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_8; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_9; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_10; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_11; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_12; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_13; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_14; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_15; // @[PRNG.scala 82:22]
  wire [29:0] MaxPeriodFibonacciLFSR_io_covSum; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_metaAssert; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_metaReset; // @[PRNG.scala 82:22]
  wire  metaArb_io_in_0_valid; // @[DCache.scala 120:23]
  wire [39:0] metaArb_io_in_0_bits_addr; // @[DCache.scala 120:23]
  wire [5:0] metaArb_io_in_0_bits_idx; // @[DCache.scala 120:23]
  wire [21:0] metaArb_io_in_0_bits_data; // @[DCache.scala 120:23]
  wire  metaArb_io_in_1_valid; // @[DCache.scala 120:23]
  wire [39:0] metaArb_io_in_1_bits_addr; // @[DCache.scala 120:23]
  wire [5:0] metaArb_io_in_1_bits_idx; // @[DCache.scala 120:23]
  wire [21:0] metaArb_io_in_1_bits_data; // @[DCache.scala 120:23]
  wire  metaArb_io_in_2_valid; // @[DCache.scala 120:23]
  wire [39:0] metaArb_io_in_2_bits_addr; // @[DCache.scala 120:23]
  wire [5:0] metaArb_io_in_2_bits_idx; // @[DCache.scala 120:23]
  wire [3:0] metaArb_io_in_2_bits_way_en; // @[DCache.scala 120:23]
  wire [21:0] metaArb_io_in_2_bits_data; // @[DCache.scala 120:23]
  wire  metaArb_io_in_3_valid; // @[DCache.scala 120:23]
  wire [39:0] metaArb_io_in_3_bits_addr; // @[DCache.scala 120:23]
  wire [5:0] metaArb_io_in_3_bits_idx; // @[DCache.scala 120:23]
  wire [3:0] metaArb_io_in_3_bits_way_en; // @[DCache.scala 120:23]
  wire [21:0] metaArb_io_in_3_bits_data; // @[DCache.scala 120:23]
  wire  metaArb_io_in_4_ready; // @[DCache.scala 120:23]
  wire  metaArb_io_in_4_valid; // @[DCache.scala 120:23]
  wire [39:0] metaArb_io_in_4_bits_addr; // @[DCache.scala 120:23]
  wire [5:0] metaArb_io_in_4_bits_idx; // @[DCache.scala 120:23]
  wire [3:0] metaArb_io_in_4_bits_way_en; // @[DCache.scala 120:23]
  wire [21:0] metaArb_io_in_4_bits_data; // @[DCache.scala 120:23]
  wire  metaArb_io_in_5_ready; // @[DCache.scala 120:23]
  wire  metaArb_io_in_5_valid; // @[DCache.scala 120:23]
  wire [39:0] metaArb_io_in_5_bits_addr; // @[DCache.scala 120:23]
  wire [5:0] metaArb_io_in_5_bits_idx; // @[DCache.scala 120:23]
  wire  metaArb_io_in_6_ready; // @[DCache.scala 120:23]
  wire  metaArb_io_in_6_valid; // @[DCache.scala 120:23]
  wire [39:0] metaArb_io_in_6_bits_addr; // @[DCache.scala 120:23]
  wire [5:0] metaArb_io_in_6_bits_idx; // @[DCache.scala 120:23]
  wire [3:0] metaArb_io_in_6_bits_way_en; // @[DCache.scala 120:23]
  wire [21:0] metaArb_io_in_6_bits_data; // @[DCache.scala 120:23]
  wire  metaArb_io_in_7_ready; // @[DCache.scala 120:23]
  wire  metaArb_io_in_7_valid; // @[DCache.scala 120:23]
  wire [39:0] metaArb_io_in_7_bits_addr; // @[DCache.scala 120:23]
  wire [5:0] metaArb_io_in_7_bits_idx; // @[DCache.scala 120:23]
  wire [3:0] metaArb_io_in_7_bits_way_en; // @[DCache.scala 120:23]
  wire [21:0] metaArb_io_in_7_bits_data; // @[DCache.scala 120:23]
  wire  metaArb_io_out_valid; // @[DCache.scala 120:23]
  wire  metaArb_io_out_bits_write; // @[DCache.scala 120:23]
  wire [39:0] metaArb_io_out_bits_addr; // @[DCache.scala 120:23]
  wire [5:0] metaArb_io_out_bits_idx; // @[DCache.scala 120:23]
  wire [3:0] metaArb_io_out_bits_way_en; // @[DCache.scala 120:23]
  wire [21:0] metaArb_io_out_bits_data; // @[DCache.scala 120:23]
  wire [29:0] metaArb_io_covSum; // @[DCache.scala 120:23]
  wire  metaArb_metaAssert; // @[DCache.scala 120:23]
  reg [21:0] tag_array_0 [0:63]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_0;
  wire [21:0] tag_array_0_s1_meta_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_0_s1_meta_addr; // @[DescribedSRAM.scala 23:26]
  wire [21:0] tag_array_0__T_260_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_0__T_260_addr; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_0__T_260_mask; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_0__T_260_en; // @[DescribedSRAM.scala 23:26]
  reg  tag_array_0_s1_meta_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] tag_array_0_s1_meta_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg [21:0] tag_array_1 [0:63]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_3;
  wire [21:0] tag_array_1_s1_meta_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_1_s1_meta_addr; // @[DescribedSRAM.scala 23:26]
  wire [21:0] tag_array_1__T_260_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_1__T_260_addr; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_1__T_260_mask; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_1__T_260_en; // @[DescribedSRAM.scala 23:26]
  reg  tag_array_1_s1_meta_en_pipe_0;
  reg [31:0] _RAND_4;
  reg [5:0] tag_array_1_s1_meta_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [21:0] tag_array_2 [0:63]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_6;
  wire [21:0] tag_array_2_s1_meta_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_2_s1_meta_addr; // @[DescribedSRAM.scala 23:26]
  wire [21:0] tag_array_2__T_260_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_2__T_260_addr; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_2__T_260_mask; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_2__T_260_en; // @[DescribedSRAM.scala 23:26]
  reg  tag_array_2_s1_meta_en_pipe_0;
  reg [31:0] _RAND_7;
  reg [5:0] tag_array_2_s1_meta_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [21:0] tag_array_3 [0:63]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_9;
  wire [21:0] tag_array_3_s1_meta_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_3_s1_meta_addr; // @[DescribedSRAM.scala 23:26]
  wire [21:0] tag_array_3__T_260_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_3__T_260_addr; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_3__T_260_mask; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_3__T_260_en; // @[DescribedSRAM.scala 23:26]
  reg  tag_array_3_s1_meta_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [5:0] tag_array_3_s1_meta_addr_pipe_0;
  reg [31:0] _RAND_11;
  wire  data_clock; // @[DCache.scala 130:20]
  wire  data_io_req_valid; // @[DCache.scala 130:20]
  wire [11:0] data_io_req_bits_addr; // @[DCache.scala 130:20]
  wire  data_io_req_bits_write; // @[DCache.scala 130:20]
  wire [63:0] data_io_req_bits_wdata; // @[DCache.scala 130:20]
  wire [7:0] data_io_req_bits_eccMask; // @[DCache.scala 130:20]
  wire [3:0] data_io_req_bits_way_en; // @[DCache.scala 130:20]
  wire [63:0] data_io_resp_0; // @[DCache.scala 130:20]
  wire [63:0] data_io_resp_1; // @[DCache.scala 130:20]
  wire [63:0] data_io_resp_2; // @[DCache.scala 130:20]
  wire [63:0] data_io_resp_3; // @[DCache.scala 130:20]
  wire [29:0] data_io_covSum; // @[DCache.scala 130:20]
  wire  data_metaAssert; // @[DCache.scala 130:20]
  wire  data_metaReset; // @[DCache.scala 130:20]
  wire  dataArb_io_in_0_valid; // @[DCache.scala 131:23]
  wire [11:0] dataArb_io_in_0_bits_addr; // @[DCache.scala 131:23]
  wire  dataArb_io_in_0_bits_write; // @[DCache.scala 131:23]
  wire [63:0] dataArb_io_in_0_bits_wdata; // @[DCache.scala 131:23]
  wire [7:0] dataArb_io_in_0_bits_eccMask; // @[DCache.scala 131:23]
  wire [3:0] dataArb_io_in_0_bits_way_en; // @[DCache.scala 131:23]
  wire  dataArb_io_in_1_ready; // @[DCache.scala 131:23]
  wire  dataArb_io_in_1_valid; // @[DCache.scala 131:23]
  wire [11:0] dataArb_io_in_1_bits_addr; // @[DCache.scala 131:23]
  wire  dataArb_io_in_1_bits_write; // @[DCache.scala 131:23]
  wire [63:0] dataArb_io_in_1_bits_wdata; // @[DCache.scala 131:23]
  wire [7:0] dataArb_io_in_1_bits_eccMask; // @[DCache.scala 131:23]
  wire [3:0] dataArb_io_in_1_bits_way_en; // @[DCache.scala 131:23]
  wire  dataArb_io_in_2_ready; // @[DCache.scala 131:23]
  wire  dataArb_io_in_2_valid; // @[DCache.scala 131:23]
  wire [11:0] dataArb_io_in_2_bits_addr; // @[DCache.scala 131:23]
  wire [63:0] dataArb_io_in_2_bits_wdata; // @[DCache.scala 131:23]
  wire [7:0] dataArb_io_in_2_bits_eccMask; // @[DCache.scala 131:23]
  wire  dataArb_io_in_3_ready; // @[DCache.scala 131:23]
  wire  dataArb_io_in_3_valid; // @[DCache.scala 131:23]
  wire [11:0] dataArb_io_in_3_bits_addr; // @[DCache.scala 131:23]
  wire [63:0] dataArb_io_in_3_bits_wdata; // @[DCache.scala 131:23]
  wire [7:0] dataArb_io_in_3_bits_eccMask; // @[DCache.scala 131:23]
  wire  dataArb_io_out_valid; // @[DCache.scala 131:23]
  wire [11:0] dataArb_io_out_bits_addr; // @[DCache.scala 131:23]
  wire  dataArb_io_out_bits_write; // @[DCache.scala 131:23]
  wire [63:0] dataArb_io_out_bits_wdata; // @[DCache.scala 131:23]
  wire [7:0] dataArb_io_out_bits_eccMask; // @[DCache.scala 131:23]
  wire [3:0] dataArb_io_out_bits_way_en; // @[DCache.scala 131:23]
  wire [29:0] dataArb_io_covSum; // @[DCache.scala 131:23]
  wire  dataArb_metaAssert; // @[DCache.scala 131:23]
  wire [7:0] amoalu_io_mask; // @[DCache.scala 881:26]
  wire [4:0] amoalu_io_cmd; // @[DCache.scala 881:26]
  wire [63:0] amoalu_io_lhs; // @[DCache.scala 881:26]
  wire [63:0] amoalu_io_rhs; // @[DCache.scala 881:26]
  wire [63:0] amoalu_io_out; // @[DCache.scala 881:26]
  wire [29:0] amoalu_io_covSum; // @[DCache.scala 881:26]
  wire  amoalu_metaAssert; // @[DCache.scala 881:26]
  wire [7:0] _T_7; // @[PRNG.scala 86:17]
  wire [15:0] _T_15; // @[PRNG.scala 86:17]
  wire  _T_16; // @[Decoupled.scala 40:37]
  reg  s1_valid; // @[DCache.scala 159:21]
  reg [31:0] _RAND_12;
  reg [2:0] blockProbeAfterGrantCount; // @[DCache.scala 611:38]
  reg [31:0] _RAND_13;
  wire  _T_2882; // @[DCache.scala 709:65]
  reg [6:0] lrscCount; // @[DCache.scala 423:22]
  reg [31:0] _RAND_14;
  wire  lrscValid; // @[DCache.scala 424:29]
  wire  block_probe_for_core_progress; // @[DCache.scala 709:69]
  reg  s1_probe; // @[DCache.scala 160:21]
  reg [31:0] _RAND_15;
  reg  s2_probe; // @[DCache.scala 285:21]
  reg [31:0] _RAND_16;
  wire  _T_381; // @[DCache.scala 286:34]
  reg [2:0] release_state; // @[DCache.scala 199:26]
  reg [31:0] _RAND_17;
  wire  _T_382; // @[DCache.scala 286:63]
  wire  releaseInFlight; // @[DCache.scala 286:46]
  reg  release_ack_wait; // @[DCache.scala 197:29]
  reg [31:0] _RAND_18;
  reg [31:0] release_ack_addr; // @[DCache.scala 198:29]
  reg [31:0] _RAND_19;
  wire [31:0] _T_2883; // @[DCache.scala 710:88]
  wire  _T_2885; // @[DCache.scala 710:124]
  wire  block_probe_for_pending_release_ack; // @[DCache.scala 710:62]
  wire  _T_2886; // @[DCache.scala 711:50]
  reg  grantInProgress; // @[DCache.scala 610:28]
  reg [31:0] _RAND_20;
  wire  block_probe_for_ordering; // @[DCache.scala 711:89]
  wire  _T_2890; // @[DCache.scala 713:79]
  wire  _T_2891; // @[DCache.scala 713:107]
  reg  s2_valid; // @[DCache.scala 283:21]
  reg [31:0] _RAND_21;
  wire  _T_2892; // @[DCache.scala 713:119]
  wire  tl_out__b_ready; // @[DCache.scala 713:44]
  wire  _T_17; // @[Decoupled.scala 40:37]
  reg [1:0] probe_bits_param; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [3:0] probe_bits_size; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg  probe_bits_source; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [31:0] probe_bits_address; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  wire  s1_valid_masked; // @[DCache.scala 163:34]
  wire  s2_meta_error; // @[DCache.scala 314:83]
  reg [1:0] s2_probe_state_state; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  wire [3:0] _T_680; // @[Cat.scala 29:58]
  wire  _T_737; // @[Misc.scala 55:20]
  wire  _T_733; // @[Misc.scala 55:20]
  wire  _T_729; // @[Misc.scala 55:20]
  wire  _T_725; // @[Misc.scala 55:20]
  wire  _T_721; // @[Misc.scala 55:20]
  wire  _T_717; // @[Misc.scala 55:20]
  wire  _T_713; // @[Misc.scala 55:20]
  wire  _T_709; // @[Misc.scala 55:20]
  wire  _T_705; // @[Misc.scala 55:20]
  wire  _T_701; // @[Misc.scala 55:20]
  wire  _T_697; // @[Misc.scala 55:20]
  wire  _T_693; // @[Misc.scala 55:20]
  wire  _T_710; // @[Misc.scala 37:9]
  wire  _T_714; // @[Misc.scala 37:9]
  wire  _T_718; // @[Misc.scala 37:9]
  wire  _T_722; // @[Misc.scala 37:9]
  wire  _T_726; // @[Misc.scala 37:9]
  wire  _T_730; // @[Misc.scala 37:9]
  wire  _T_734; // @[Misc.scala 37:9]
  wire  s2_prb_ack_data; // @[Misc.scala 37:9]
  wire  _T_2943; // @[Metadata.scala 50:45]
  reg [8:0] _T_2906; // @[Edges.scala 230:27]
  reg [31:0] _RAND_27;
  wire  _T_2909; // @[Edges.scala 233:25]
  wire  _T_2954; // @[package.scala 15:47]
  wire  _T_2955; // @[package.scala 15:47]
  wire  _T_2956; // @[package.scala 64:59]
  wire  _T_2953; // @[DCache.scala 779:25]
  wire  _T_2952; // @[DCache.scala 774:25]
  wire [2:0] _GEN_314; // @[DCache.scala 779:48]
  wire [2:0] tl_out__c_bits_opcode; // @[DCache.scala 783:81]
  wire [3:0] tl_out__c_bits_size; // @[DCache.scala 783:81]
  wire [26:0] _T_2900; // @[package.scala 212:77]
  wire [8:0] _T_2903; // @[Edges.scala 221:59]
  wire [8:0] _T_2905; // @[Edges.scala 222:14]
  wire  _T_2910; // @[Edges.scala 233:47]
  wire  c_last; // @[Edges.scala 233:37]
  wire  _T_2951; // @[DCache.scala 770:25]
  reg  s2_release_data_valid; // @[DCache.scala 724:34]
  reg [31:0] _RAND_28;
  wire  c_first; // @[Edges.scala 232:25]
  wire  _T_2925; // @[DCache.scala 732:56]
  wire  _T_2927; // @[DCache.scala 732:43]
  wire  _GEN_263; // @[DCache.scala 748:36]
  wire  _GEN_273; // @[DCache.scala 746:28]
  wire  _GEN_284; // @[DCache.scala 744:21]
  wire  _GEN_301; // @[DCache.scala 770:47]
  wire  tl_out__c_valid; // @[DCache.scala 774:48]
  wire  _T_2898; // @[Decoupled.scala 40:37]
  wire  releaseDone; // @[Edges.scala 234:22]
  wire  _GEN_261; // @[DCache.scala 750:45]
  wire  _GEN_271; // @[DCache.scala 748:36]
  wire  probeNack; // @[DCache.scala 746:28]
  reg [4:0] s1_req_cmd; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  wire  _T_30; // @[Consts.scala 82:31]
  wire  _T_31; // @[Consts.scala 82:48]
  wire  _T_32; // @[Consts.scala 82:41]
  wire  _T_33; // @[Consts.scala 82:65]
  wire  _T_34; // @[Consts.scala 82:58]
  wire  _T_35; // @[package.scala 15:47]
  wire  _T_36; // @[package.scala 15:47]
  wire  _T_39; // @[package.scala 64:59]
  wire  _T_37; // @[package.scala 15:47]
  wire  _T_40; // @[package.scala 64:59]
  wire  _T_38; // @[package.scala 15:47]
  wire  _T_41; // @[package.scala 64:59]
  wire  _T_42; // @[package.scala 15:47]
  wire  _T_43; // @[package.scala 15:47]
  wire  _T_47; // @[package.scala 64:59]
  wire  _T_44; // @[package.scala 15:47]
  wire  _T_48; // @[package.scala 64:59]
  wire  _T_45; // @[package.scala 15:47]
  wire  _T_49; // @[package.scala 64:59]
  wire  _T_46; // @[package.scala 15:47]
  wire  _T_50; // @[package.scala 64:59]
  wire  _T_51; // @[Consts.scala 80:44]
  wire  s1_read; // @[Consts.scala 82:75]
  reg [4:0] s2_req_cmd; // @[DCache.scala 291:19]
  reg [31:0] _RAND_30;
  wire  _T_418; // @[Consts.scala 83:32]
  wire  _T_419; // @[Consts.scala 83:49]
  wire  _T_420; // @[Consts.scala 83:42]
  wire  _T_421; // @[Consts.scala 83:66]
  wire  _T_422; // @[Consts.scala 83:59]
  wire  _T_423; // @[package.scala 15:47]
  wire  _T_424; // @[package.scala 15:47]
  wire  _T_427; // @[package.scala 64:59]
  wire  _T_425; // @[package.scala 15:47]
  wire  _T_428; // @[package.scala 64:59]
  wire  _T_426; // @[package.scala 15:47]
  wire  _T_429; // @[package.scala 64:59]
  wire  _T_430; // @[package.scala 15:47]
  wire  _T_431; // @[package.scala 15:47]
  wire  _T_435; // @[package.scala 64:59]
  wire  _T_432; // @[package.scala 15:47]
  wire  _T_436; // @[package.scala 64:59]
  wire  _T_433; // @[package.scala 15:47]
  wire  _T_437; // @[package.scala 64:59]
  wire  _T_434; // @[package.scala 15:47]
  wire  _T_438; // @[package.scala 64:59]
  wire  _T_439; // @[Consts.scala 80:44]
  wire  s2_write; // @[Consts.scala 83:76]
  wire  _T_1017; // @[DCache.scala 456:39]
  reg  pstore1_held; // @[DCache.scala 455:25]
  reg [31:0] _RAND_31;
  wire  pstore1_valid_likely; // @[DCache.scala 456:51]
  reg [39:0] pstore1_addr; // @[Reg.scala 15:16]
  reg [63:0] _RAND_32;
  reg [39:0] s1_req_addr; // @[Reg.scala 15:16]
  reg [63:0] _RAND_33;
  wire  _T_1178; // @[DCache.scala 508:31]
  wire  _T_52; // @[Consts.scala 83:32]
  wire  _T_53; // @[Consts.scala 83:49]
  wire  _T_54; // @[Consts.scala 83:42]
  wire  _T_56; // @[Consts.scala 83:59]
  wire  s1_write; // @[Consts.scala 83:76]
  reg [7:0] pstore1_mask; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  wire  _T_1194; // @[DCache.scala 1076:66]
  wire  _T_1193; // @[DCache.scala 1076:66]
  wire  _T_1192; // @[DCache.scala 1076:66]
  wire  _T_1191; // @[DCache.scala 1076:66]
  wire  _T_1190; // @[DCache.scala 1076:66]
  wire  _T_1189; // @[DCache.scala 1076:66]
  wire  _T_1188; // @[DCache.scala 1076:66]
  wire  _T_1187; // @[DCache.scala 1076:66]
  wire [7:0] _T_1201; // @[Cat.scala 29:58]
  wire [7:0] _T_1216; // @[Cat.scala 29:58]
  reg [1:0] s1_req_size; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  wire  _T_340; // @[AMOALU.scala 17:57]
  wire  _T_342; // @[AMOALU.scala 17:46]
  wire  _T_344; // @[AMOALU.scala 18:22]
  wire [1:0] _T_345; // @[Cat.scala 29:58]
  wire [1:0] _T_347; // @[AMOALU.scala 17:22]
  wire  _T_348; // @[AMOALU.scala 17:57]
  wire [1:0] _T_349; // @[AMOALU.scala 17:51]
  wire [1:0] _T_350; // @[AMOALU.scala 17:46]
  wire [1:0] _T_352; // @[AMOALU.scala 18:22]
  wire [3:0] _T_353; // @[Cat.scala 29:58]
  wire [3:0] _T_355; // @[AMOALU.scala 17:22]
  wire  _T_356; // @[AMOALU.scala 17:57]
  wire [3:0] _T_357; // @[AMOALU.scala 17:51]
  wire [3:0] _T_358; // @[AMOALU.scala 17:46]
  wire [3:0] _T_360; // @[AMOALU.scala 18:22]
  wire [7:0] s1_mask_xwr; // @[Cat.scala 29:58]
  wire  _T_1232; // @[DCache.scala 1076:66]
  wire  _T_1231; // @[DCache.scala 1076:66]
  wire  _T_1230; // @[DCache.scala 1076:66]
  wire  _T_1229; // @[DCache.scala 1076:66]
  wire  _T_1228; // @[DCache.scala 1076:66]
  wire  _T_1227; // @[DCache.scala 1076:66]
  wire  _T_1226; // @[DCache.scala 1076:66]
  wire  _T_1225; // @[DCache.scala 1076:66]
  wire [7:0] _T_1239; // @[Cat.scala 29:58]
  wire [7:0] _T_1254; // @[Cat.scala 29:58]
  wire [7:0] _T_1255; // @[DCache.scala 509:38]
  wire  _T_1256; // @[DCache.scala 509:66]
  wire [7:0] _T_1257; // @[DCache.scala 509:77]
  wire  _T_1258; // @[DCache.scala 509:92]
  wire  _T_1259; // @[DCache.scala 509:8]
  wire  _T_1260; // @[DCache.scala 508:68]
  wire  _T_1261; // @[DCache.scala 511:27]
  reg  pstore2_valid; // @[DCache.scala 452:26]
  reg [31:0] _RAND_36;
  reg [39:0] pstore2_addr; // @[Reg.scala 15:16]
  reg [63:0] _RAND_37;
  wire  _T_1264; // @[DCache.scala 508:31]
  reg [7:0] mask; // @[DCache.scala 482:19]
  reg [31:0] _RAND_38;
  wire  _T_1280; // @[DCache.scala 1076:66]
  wire  _T_1279; // @[DCache.scala 1076:66]
  wire  _T_1278; // @[DCache.scala 1076:66]
  wire  _T_1277; // @[DCache.scala 1076:66]
  wire  _T_1276; // @[DCache.scala 1076:66]
  wire  _T_1275; // @[DCache.scala 1076:66]
  wire  _T_1274; // @[DCache.scala 1076:66]
  wire  _T_1273; // @[DCache.scala 1076:66]
  wire [7:0] _T_1287; // @[Cat.scala 29:58]
  wire [7:0] _T_1302; // @[Cat.scala 29:58]
  wire [7:0] _T_1341; // @[DCache.scala 509:38]
  wire  _T_1342; // @[DCache.scala 509:66]
  wire [7:0] _T_1343; // @[DCache.scala 509:77]
  wire  _T_1344; // @[DCache.scala 509:92]
  wire  _T_1345; // @[DCache.scala 509:8]
  wire  _T_1346; // @[DCache.scala 508:68]
  wire  _T_1347; // @[DCache.scala 512:21]
  wire  s1_hazard; // @[DCache.scala 511:69]
  wire  s1_raw_hazard; // @[DCache.scala 513:31]
  wire  _T_1348; // @[DCache.scala 518:18]
  wire [5:0] _T_378; // @[DCache.scala 284:54]
  wire  _T_379; // @[DCache.scala 284:61]
  wire  s2_valid_no_xcpt; // @[DCache.scala 284:35]
  reg  s2_not_nacked_in_s1; // @[DCache.scala 287:36]
  reg [31:0] _RAND_39;
  wire  s2_valid_masked; // @[DCache.scala 289:42]
  wire  _T_644; // @[DCache.scala 349:71]
  wire  _T_539; // @[Consts.scala 84:54]
  wire  _T_540; // @[Consts.scala 84:47]
  wire  _T_541; // @[Consts.scala 84:71]
  wire  _T_542; // @[Consts.scala 84:64]
  reg [1:0] s2_hit_state_state; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  wire [3:0] _T_544; // @[Cat.scala 29:58]
  wire  _T_602; // @[Misc.scala 48:20]
  wire  _T_599; // @[Misc.scala 48:20]
  wire  _T_596; // @[Misc.scala 48:20]
  wire  _T_593; // @[Misc.scala 48:20]
  wire  _T_590; // @[Misc.scala 48:20]
  wire  _T_587; // @[Misc.scala 48:20]
  wire  _T_584; // @[Misc.scala 48:20]
  wire  _T_581; // @[Misc.scala 48:20]
  wire  _T_578; // @[Misc.scala 48:20]
  wire  _T_575; // @[Misc.scala 48:20]
  wire  _T_572; // @[Misc.scala 48:20]
  wire  _T_569; // @[Misc.scala 48:20]
  wire  _T_588; // @[Misc.scala 34:9]
  wire  _T_591; // @[Misc.scala 34:9]
  wire  _T_594; // @[Misc.scala 34:9]
  wire  _T_597; // @[Misc.scala 34:9]
  wire  _T_600; // @[Misc.scala 34:9]
  wire  s2_hit; // @[Misc.scala 34:9]
  wire  s2_valid_hit_maybe_flush_pre_data_ecc_and_waw; // @[DCache.scala 349:89]
  wire  _T_396; // @[Consts.scala 82:31]
  wire  _T_398; // @[Consts.scala 82:41]
  wire  _T_400; // @[Consts.scala 82:58]
  wire  s2_read; // @[Consts.scala 82:75]
  wire  s2_readwrite; // @[DCache.scala 306:30]
  wire  s2_valid_hit_pre_data_ecc_and_waw; // @[DCache.scala 370:89]
  wire [1:0] _T_571; // @[Misc.scala 34:36]
  wire [1:0] _T_574; // @[Misc.scala 34:36]
  wire [1:0] _T_577; // @[Misc.scala 34:36]
  wire [1:0] _T_580; // @[Misc.scala 34:36]
  wire [1:0] _T_583; // @[Misc.scala 34:36]
  wire [1:0] _T_586; // @[Misc.scala 34:36]
  wire [1:0] _T_589; // @[Misc.scala 34:36]
  wire [1:0] _T_592; // @[Misc.scala 34:36]
  wire [1:0] _T_595; // @[Misc.scala 34:36]
  wire [1:0] _T_598; // @[Misc.scala 34:36]
  wire [1:0] _T_601; // @[Misc.scala 34:36]
  wire [1:0] s2_grow_param; // @[Misc.scala 34:36]
  wire  _T_804; // @[Metadata.scala 46:46]
  wire  s2_update_meta; // @[Metadata.scala 47:40]
  wire  _T_823; // @[DCache.scala 397:62]
  wire  _T_824; // @[DCache.scala 397:24]
  wire  s1_readwrite; // @[DCache.scala 185:30]
  wire  _T_74; // @[DCache.scala 187:34]
  wire  s1_flush_line; // @[DCache.scala 187:50]
  wire  _T_227; // @[DCache.scala 229:38]
  wire  _T_228; // @[DCache.scala 229:69]
  wire  s1_cmd_uses_tlb; // @[DCache.scala 229:55]
  wire  _T_242; // @[DCache.scala 235:39]
  wire  _T_243; // @[DCache.scala 235:58]
  wire  _GEN_118; // @[DCache.scala 397:82]
  wire  _GEN_142; // @[DCache.scala 518:36]
  wire  _GEN_282; // @[DCache.scala 759:24]
  wire  s1_nack; // @[DCache.scala 744:21]
  wire  s1_valid_not_nacked; // @[DCache.scala 164:38]
  wire  s0_clk_en; // @[DCache.scala 167:40]
  wire [39:0] s0_req_addr; // @[Cat.scala 29:58]
  wire  s0_req_phys; // @[DCache.scala 171:34]
  reg [6:0] s1_req_tag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg  s1_req_signed; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [39:0] s1_tlb_req_vaddr; // @[Reg.scala 15:16]
  reg [63:0] _RAND_43;
  reg  s1_tlb_req_passthrough; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [1:0] s1_tlb_req_size; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [4:0] s1_tlb_req_cmd; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  wire  s1_sfence; // @[DCache.scala 186:30]
  reg  s1_flush_valid; // @[DCache.scala 188:27]
  reg [31:0] _RAND_47;
  reg  cached_grant_wait; // @[DCache.scala 196:30]
  reg [31:0] _RAND_48;
  wire  inWriteback; // @[package.scala 64:59]
  wire  _T_78; // @[DCache.scala 203:38]
  wire  _T_80; // @[DCache.scala 203:51]
  wire  _T_82; // @[DCache.scala 203:73]
  reg  uncachedInFlight_0; // @[DCache.scala 206:33]
  reg [31:0] _RAND_49;
  reg [39:0] uncachedReqs_0_addr; // @[DCache.scala 207:25]
  reg [63:0] _RAND_50;
  reg [6:0] uncachedReqs_0_tag; // @[DCache.scala 207:25]
  reg [31:0] _RAND_51;
  reg [1:0] uncachedReqs_0_size; // @[DCache.scala 207:25]
  reg [31:0] _RAND_52;
  reg  uncachedReqs_0_signed; // @[DCache.scala 207:25]
  reg [31:0] _RAND_53;
  wire  _T_84; // @[Consts.scala 82:31]
  wire  _T_85; // @[Consts.scala 82:48]
  wire  _T_86; // @[Consts.scala 82:41]
  wire  _T_87; // @[Consts.scala 82:65]
  wire  _T_88; // @[Consts.scala 82:58]
  wire  _T_89; // @[package.scala 15:47]
  wire  _T_90; // @[package.scala 15:47]
  wire  _T_91; // @[package.scala 15:47]
  wire  _T_92; // @[package.scala 15:47]
  wire  _T_93; // @[package.scala 64:59]
  wire  _T_94; // @[package.scala 64:59]
  wire  _T_95; // @[package.scala 64:59]
  wire  _T_96; // @[package.scala 15:47]
  wire  _T_97; // @[package.scala 15:47]
  wire  _T_98; // @[package.scala 15:47]
  wire  _T_99; // @[package.scala 15:47]
  wire  _T_100; // @[package.scala 15:47]
  wire  _T_101; // @[package.scala 64:59]
  wire  _T_102; // @[package.scala 64:59]
  wire  _T_103; // @[package.scala 64:59]
  wire  _T_104; // @[package.scala 64:59]
  wire  _T_105; // @[Consts.scala 80:44]
  wire  s0_read; // @[Consts.scala 82:75]
  wire  _T_106; // @[package.scala 15:47]
  wire  _T_107; // @[package.scala 15:47]
  wire  _T_108; // @[package.scala 64:59]
  wire  res; // @[DCache.scala 1080:15]
  wire  _T_135; // @[Consts.scala 83:49]
  wire  _T_136; // @[Consts.scala 83:42]
  wire  _T_138; // @[Consts.scala 83:59]
  wire  _T_156; // @[Consts.scala 83:76]
  wire  _T_160; // @[DCache.scala 1086:23]
  wire  _T_161; // @[DCache.scala 1085:21]
  wire  _T_163; // @[DCache.scala 1081:28]
  wire  _T_165; // @[DCache.scala 1081:11]
  wire  _T_167; // @[DCache.scala 212:46]
  wire  _T_171; // @[DCache.scala 218:33]
  wire  _GEN_28; // @[DCache.scala 218:45]
  wire  _T_223; // @[DCache.scala 219:75]
  wire  _T_224; // @[DCache.scala 219:54]
  reg  s1_did_read; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  wire  _GEN_30; // @[DCache.scala 226:34]
  wire  _T_237; // @[DCache.scala 234:27]
  wire  _T_239; // @[DCache.scala 234:53]
  wire  _GEN_31; // @[DCache.scala 234:79]
  wire [31:0] s1_paddr; // @[Cat.scala 29:58]
  wire [1:0] s1_victim_way; // @[package.scala 143:13]
  wire [21:0] _T_266;
  wire [19:0] s1_meta_uncorrected_0_tag; // @[DCache.scala 267:80]
  wire [1:0] s1_meta_uncorrected_0_coh_state; // @[DCache.scala 267:80]
  wire [21:0] _T_269;
  wire [19:0] s1_meta_uncorrected_1_tag; // @[DCache.scala 267:80]
  wire [1:0] s1_meta_uncorrected_1_coh_state; // @[DCache.scala 267:80]
  wire [21:0] _T_272;
  wire [19:0] s1_meta_uncorrected_2_tag; // @[DCache.scala 267:80]
  wire [1:0] s1_meta_uncorrected_2_coh_state; // @[DCache.scala 267:80]
  wire [21:0] _T_275;
  wire [19:0] s1_meta_uncorrected_3_tag; // @[DCache.scala 267:80]
  wire [1:0] s1_meta_uncorrected_3_coh_state; // @[DCache.scala 267:80]
  wire [19:0] s1_tag; // @[DCache.scala 268:29]
  wire  _T_278; // @[Metadata.scala 50:45]
  wire  _T_279; // @[DCache.scala 269:83]
  wire  _T_280; // @[DCache.scala 269:74]
  wire  _T_281; // @[Metadata.scala 50:45]
  wire  _T_282; // @[DCache.scala 269:83]
  wire  _T_283; // @[DCache.scala 269:74]
  wire  _T_284; // @[Metadata.scala 50:45]
  wire  _T_285; // @[DCache.scala 269:83]
  wire  _T_286; // @[DCache.scala 269:74]
  wire  _T_287; // @[Metadata.scala 50:45]
  wire  _T_288; // @[DCache.scala 269:83]
  wire  _T_289; // @[DCache.scala 269:74]
  wire [3:0] s1_meta_hit_way; // @[Cat.scala 29:58]
  wire  _T_295; // @[DCache.scala 271:59]
  wire [1:0] _T_296; // @[DCache.scala 271:41]
  wire  _T_299; // @[DCache.scala 271:59]
  wire [1:0] _T_300; // @[DCache.scala 271:41]
  wire  _T_303; // @[DCache.scala 271:59]
  wire [1:0] _T_304; // @[DCache.scala 271:41]
  wire  _T_307; // @[DCache.scala 271:59]
  wire [1:0] _T_308; // @[DCache.scala 271:41]
  wire [1:0] _T_309; // @[DCache.scala 272:19]
  wire [1:0] _T_310; // @[DCache.scala 272:19]
  wire [1:0] s1_meta_hit_state_state; // @[DCache.scala 272:19]
  wire  _T_316; // @[package.scala 32:86]
  wire  _T_318; // @[package.scala 32:86]
  wire  _T_320; // @[package.scala 32:86]
  wire  s2_hit_valid; // @[Metadata.scala 50:45]
  reg [3:0] s2_hit_way; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [1:0] _T_672; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  wire [3:0] _T_673; // @[OneHot.scala 58:35]
  wire [3:0] s2_victim_way; // @[DCache.scala 383:26]
  reg [3:0] s2_probe_way; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  wire [3:0] releaseWay; // @[DCache.scala 783:81]
  wire [3:0] _T_321; // @[DCache.scala 275:61]
  wire [31:0] _T_332; // @[Cat.scala 29:58]
  wire [31:0] _T_335; // @[Cat.scala 29:58]
  wire [63:0] _T_336; // @[Cat.scala 29:58]
  wire  _T_363; // @[DCache.scala 281:28]
  wire  _T_367; // @[DCache.scala 281:93]
  wire  _T_368; // @[DCache.scala 281:53]
  wire  _T_370; // @[DCache.scala 281:9]
  wire  _T_373; // @[DCache.scala 283:43]
  reg [39:0] s2_req_addr; // @[DCache.scala 291:19]
  reg [63:0] _RAND_58;
  reg [6:0] s2_req_tag; // @[DCache.scala 291:19]
  reg [31:0] _RAND_59;
  reg [1:0] s2_req_size; // @[DCache.scala 291:19]
  reg [31:0] _RAND_60;
  reg  s2_req_signed; // @[DCache.scala 291:19]
  reg [31:0] _RAND_61;
  wire  _T_385; // @[DCache.scala 292:37]
  wire  s2_cmd_flush_line; // @[DCache.scala 293:54]
  reg  s2_tlb_xcpt_pf_ld; // @[DCache.scala 294:24]
  reg [31:0] _RAND_62;
  reg  s2_tlb_xcpt_pf_st; // @[DCache.scala 294:24]
  reg [31:0] _RAND_63;
  reg  s2_tlb_xcpt_ae_ld; // @[DCache.scala 294:24]
  reg [31:0] _RAND_64;
  reg  s2_tlb_xcpt_ae_st; // @[DCache.scala 294:24]
  reg [31:0] _RAND_65;
  reg  s2_tlb_xcpt_ma_ld; // @[DCache.scala 294:24]
  reg [31:0] _RAND_66;
  reg  s2_tlb_xcpt_ma_st; // @[DCache.scala 294:24]
  reg [31:0] _RAND_67;
  reg  s2_pma_cacheable; // @[DCache.scala 295:19]
  reg [31:0] _RAND_68;
  wire  _T_390; // @[DCache.scala 297:29]
  wire  _T_391_cacheable; // @[DCache.scala 301:18]
  reg [39:0] _T_393; // @[Reg.scala 15:16]
  reg [63:0] _RAND_69;
  wire [39:0] s2_vaddr; // @[Cat.scala 29:58]
  reg  s2_flush_valid_pre_tag_ecc; // @[DCache.scala 307:43]
  reg [31:0] _RAND_70;
  wire  s1_meta_clk_en; // @[DCache.scala 309:62]
  reg [21:0] _T_465; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  wire [19:0] s2_meta_corrected_3_tag; // @[DCache.scala 313:99]
  wire [1:0] s2_meta_corrected_3_coh_state; // @[DCache.scala 313:99]
  wire  s2_flush_valid; // @[DCache.scala 315:51]
  wire  _T_471; // @[DCache.scala 318:23]
  wire  en; // @[DCache.scala 318:38]
  wire  _T_473; // @[DCache.scala 319:63]
  wire  word_en; // @[DCache.scala 319:22]
  wire [63:0] s1_all_data_ways_0; // @[DCache.scala 277:29 DCache.scala 277:29]
  wire [63:0] s1_all_data_ways_1; // @[DCache.scala 277:29 DCache.scala 277:29]
  wire [63:0] s1_all_data_ways_2; // @[DCache.scala 277:29 DCache.scala 277:29]
  wire [63:0] s1_all_data_ways_3; // @[DCache.scala 277:29 DCache.scala 277:29]
  wire  s1_word_en; // @[DCache.scala 329:27]
  wire  grantIsUncachedData; // @[package.scala 15:47]
  reg  blockUncachedGrant; // @[DCache.scala 693:33]
  reg [31:0] _RAND_72;
  wire  _T_2877; // @[DCache.scala 695:54]
  wire  _T_2878; // @[DCache.scala 695:31]
  wire  grantIsRefill; // @[DCache.scala 609:29]
  wire  _T_2792; // @[DCache.scala 665:23]
  wire  _T_2745; // @[package.scala 15:47]
  wire  grantIsCached; // @[package.scala 64:59]
  reg [8:0] _T_2713; // @[Edges.scala 230:27]
  reg [31:0] _RAND_73;
  wire  d_first; // @[Edges.scala 232:25]
  wire  _T_2754; // @[DCache.scala 614:50]
  wire  canAcceptCachedGrant; // @[DCache.scala 613:30]
  wire  _T_2755; // @[DCache.scala 614:69]
  wire  _T_2756; // @[DCache.scala 614:24]
  wire  _GEN_232; // @[DCache.scala 665:51]
  wire  tl_out__d_ready; // @[DCache.scala 695:68]
  wire  _T_2761; // @[Decoupled.scala 40:37]
  wire  _T_2722; // @[package.scala 15:47]
  wire  _T_2724; // @[package.scala 64:59]
  wire  _T_2723; // @[package.scala 15:47]
  wire  grantIsUncached; // @[package.scala 64:59]
  wire [4:0] _GEN_188; // @[DCache.scala 634:34]
  wire [4:0] _GEN_197; // @[DCache.scala 627:35]
  wire [4:0] _GEN_210; // @[DCache.scala 618:26]
  wire [4:0] s1_data_way; // @[DCache.scala 617:26]
  wire [4:0] _T_476; // @[DCache.scala 331:28]
  wire [63:0] _T_482; // @[Mux.scala 27:72]
  wire [63:0] _T_483; // @[Mux.scala 27:72]
  wire [63:0] _T_484; // @[Mux.scala 27:72]
  wire [63:0] _T_485; // @[Mux.scala 27:72]
  wire [63:0] _T_486; // @[Mux.scala 27:72]
  wire [63:0] _T_487; // @[Mux.scala 27:72]
  wire [63:0] _T_488; // @[Mux.scala 27:72]
  wire [63:0] _T_489; // @[Mux.scala 27:72]
  wire [63:0] _T_490; // @[Mux.scala 27:72]
  reg [63:0] s2_data; // @[Reg.scala 15:16]
  reg [63:0] _RAND_74;
  wire [31:0] _T_633; // @[Cat.scala 29:58]
  wire [31:0] _T_636; // @[Cat.scala 29:58]
  wire [63:0] s2_data_corrected; // @[Cat.scala 29:58]
  wire  s2_valid_flush_line; // @[DCache.scala 371:75]
  wire  _T_650; // @[DCache.scala 375:39]
  wire  _T_652; // @[DCache.scala 375:55]
  wire  s2_valid_miss; // @[DCache.scala 375:73]
  wire  s2_uncached; // @[DCache.scala 376:21]
  wire  _T_660; // @[DCache.scala 377:44]
  wire  _T_661; // @[DCache.scala 377:88]
  wire  s2_valid_cached_miss; // @[DCache.scala 377:60]
  wire  _T_663; // @[DCache.scala 379:79]
  wire  s2_want_victimize; // @[DCache.scala 379:125]
  wire  _T_668; // @[DCache.scala 382:49]
  wire  _T_669; // @[DCache.scala 382:92]
  wire  s2_valid_uncached_pending; // @[DCache.scala 382:64]
  reg [19:0] _T_677; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  wire [19:0] s2_victim_tag; // @[DCache.scala 384:26]
  reg [1:0] _T_679_state; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  wire [1:0] s2_victim_state_state; // @[DCache.scala 385:28]
  wire [2:0] _T_695; // @[Misc.scala 37:36]
  wire [2:0] _T_699; // @[Misc.scala 37:36]
  wire [2:0] _T_703; // @[Misc.scala 37:36]
  wire [2:0] _T_707; // @[Misc.scala 37:36]
  wire [2:0] _T_711; // @[Misc.scala 37:36]
  wire [2:0] _T_715; // @[Misc.scala 37:36]
  wire [1:0] _T_716; // @[Misc.scala 37:63]
  wire [2:0] _T_719; // @[Misc.scala 37:36]
  wire [1:0] _T_720; // @[Misc.scala 37:63]
  wire [2:0] _T_723; // @[Misc.scala 37:36]
  wire [1:0] _T_724; // @[Misc.scala 37:63]
  wire [2:0] _T_727; // @[Misc.scala 37:36]
  wire [1:0] _T_728; // @[Misc.scala 37:63]
  wire [2:0] _T_731; // @[Misc.scala 37:36]
  wire [1:0] _T_732; // @[Misc.scala 37:63]
  wire [2:0] _T_735; // @[Misc.scala 37:36]
  wire [1:0] _T_736; // @[Misc.scala 37:63]
  wire [2:0] s2_report_param; // @[Misc.scala 37:36]
  wire [1:0] probeNewCoh_state; // @[Misc.scala 37:63]
  wire [3:0] _T_745; // @[Cat.scala 29:58]
  wire  _T_758; // @[Misc.scala 55:20]
  wire [2:0] _T_760; // @[Misc.scala 37:36]
  wire  _T_762; // @[Misc.scala 55:20]
  wire [2:0] _T_764; // @[Misc.scala 37:36]
  wire  _T_766; // @[Misc.scala 55:20]
  wire [2:0] _T_768; // @[Misc.scala 37:36]
  wire  _T_770; // @[Misc.scala 55:20]
  wire [2:0] _T_772; // @[Misc.scala 37:36]
  wire  _T_774; // @[Misc.scala 55:20]
  wire  _T_775; // @[Misc.scala 37:9]
  wire [2:0] _T_776; // @[Misc.scala 37:36]
  wire  _T_778; // @[Misc.scala 55:20]
  wire  _T_779; // @[Misc.scala 37:9]
  wire [2:0] _T_780; // @[Misc.scala 37:36]
  wire [1:0] _T_781; // @[Misc.scala 37:63]
  wire  _T_782; // @[Misc.scala 55:20]
  wire  _T_783; // @[Misc.scala 37:9]
  wire [2:0] _T_784; // @[Misc.scala 37:36]
  wire [1:0] _T_785; // @[Misc.scala 37:63]
  wire  _T_786; // @[Misc.scala 55:20]
  wire  _T_787; // @[Misc.scala 37:9]
  wire [2:0] _T_788; // @[Misc.scala 37:36]
  wire [1:0] _T_789; // @[Misc.scala 37:63]
  wire  _T_790; // @[Misc.scala 55:20]
  wire  _T_791; // @[Misc.scala 37:9]
  wire [2:0] _T_792; // @[Misc.scala 37:36]
  wire [1:0] _T_793; // @[Misc.scala 37:63]
  wire  _T_794; // @[Misc.scala 55:20]
  wire  _T_795; // @[Misc.scala 37:9]
  wire [2:0] _T_796; // @[Misc.scala 37:36]
  wire [1:0] _T_797; // @[Misc.scala 37:63]
  wire  _T_798; // @[Misc.scala 55:20]
  wire  _T_799; // @[Misc.scala 37:9]
  wire [2:0] _T_800; // @[Misc.scala 37:36]
  wire [1:0] _T_801; // @[Misc.scala 37:63]
  wire  _T_802; // @[Misc.scala 55:20]
  wire  s2_victim_dirty; // @[Misc.scala 37:9]
  wire [2:0] s2_shrink_param; // @[Misc.scala 37:36]
  wire [1:0] voluntaryNewCoh_state; // @[Misc.scala 37:63]
  wire  s2_dont_nack_uncached; // @[DCache.scala 391:57]
  wire  _T_815; // @[DCache.scala 395:17]
  wire  s2_dont_nack_misc; // @[DCache.scala 392:61]
  wire  _T_818; // @[DCache.scala 396:38]
  wire  _T_820; // @[DCache.scala 396:64]
  wire  _T_831; // @[DCache.scala 401:63]
  wire  _T_832; // @[DCache.scala 401:93]
  wire [11:0] _T_848; // @[DCache.scala 405:98]
  wire [1:0] new_meta_coh_state; // @[DCache.scala 408:40]
  wire  _T_863; // @[DCache.scala 425:34]
  wire  lrscBackingOff; // @[DCache.scala 425:38]
  reg [33:0] lrscAddr; // @[DCache.scala 426:21]
  reg [63:0] _RAND_77;
  wire  lrscAddrMatch; // @[DCache.scala 427:32]
  wire  _T_866; // @[DCache.scala 428:41]
  wire  s2_sc_fail; // @[DCache.scala 428:26]
  wire  _T_868; // @[DCache.scala 429:23]
  wire  _T_870; // @[DCache.scala 429:32]
  wire  _T_871; // @[DCache.scala 429:54]
  wire [6:0] _T_878; // @[DCache.scala 433:49]
  wire  _T_879; // @[DCache.scala 434:29]
  wire  _T_887; // @[DCache.scala 443:63]
  reg [4:0] pstore1_cmd; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [63:0] pstore1_data; // @[Reg.scala 15:16]
  reg [63:0] _RAND_79;
  reg [3:0] pstore1_way; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  wire  _T_941; // @[DCache.scala 1086:23]
  wire  _T_942; // @[DCache.scala 1085:21]
  reg  pstore1_rmw; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  wire  _T_946; // @[DCache.scala 441:46]
  wire  _T_948; // @[DCache.scala 441:58]
  wire  pstore_drain_opportunistic; // @[DCache.scala 453:36]
  reg  _T_1016; // @[DCache.scala 454:56]
  reg [31:0] _RAND_82;
  wire  pstore_drain_on_miss; // @[DCache.scala 454:46]
  wire  pstore1_valid; // @[DCache.scala 458:38]
  wire  _T_1024; // @[DCache.scala 460:54]
  wire  _T_1025; // @[DCache.scala 460:85]
  wire  _T_1026; // @[DCache.scala 460:98]
  wire  pstore_drain_structural; // @[DCache.scala 460:71]
  wire  _T_1030; // @[DCache.scala 457:96]
  wire  _T_1031; // @[DCache.scala 461:63]
  wire  _T_1032; // @[DCache.scala 461:22]
  wire  _T_1034; // @[DCache.scala 461:9]
  wire  _T_1045; // @[DCache.scala 469:41]
  wire  _T_1046; // @[DCache.scala 469:58]
  wire  _T_1047; // @[DCache.scala 469:107]
  wire  _T_1048; // @[DCache.scala 469:76]
  wire  pstore_drain; // @[DCache.scala 468:48]
  wire  _T_1058; // @[DCache.scala 472:71]
  wire  _T_1062; // @[DCache.scala 473:79]
  wire  advance_pstore1; // @[DCache.scala 473:61]
  wire  _T_1064; // @[DCache.scala 474:34]
  reg [3:0] pstore2_way; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  wire [63:0] pstore1_storegen_data; // @[DCache.scala 888:27]
  reg [7:0] _T_1072; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [7:0] _T_1077; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [7:0] _T_1082; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [7:0] _T_1087; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [7:0] _T_1092; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [7:0] _T_1097; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [7:0] _T_1102; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [7:0] _T_1107; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  wire [63:0] pstore2_storegen_data; // @[Cat.scala 29:58]
  wire [39:0] _T_1132; // @[DCache.scala 500:36]
  wire [63:0] _T_1134; // @[DCache.scala 502:63]
  wire [31:0] _T_1145; // @[Cat.scala 29:58]
  wire [31:0] _T_1148; // @[Cat.scala 29:58]
  wire [7:0] _T_1152; // @[DCache.scala 504:47]
  wire  _T_1161; // @[DCache.scala 1076:66]
  wire  _T_1162; // @[DCache.scala 1076:66]
  wire  _T_1163; // @[DCache.scala 1076:66]
  wire  _T_1164; // @[DCache.scala 1076:66]
  wire  _T_1165; // @[DCache.scala 1076:66]
  wire  _T_1166; // @[DCache.scala 1076:66]
  wire  _T_1167; // @[DCache.scala 1076:66]
  wire  _T_1168; // @[DCache.scala 1076:66]
  wire [3:0] _T_1171; // @[Cat.scala 29:58]
  wire [3:0] _T_1174; // @[Cat.scala 29:58]
  wire [1:0] _T_1355; // @[DCache.scala 524:59]
  wire  a_source; // @[Mux.scala 47:69]
  wire [39:0] acquire_address; // @[DCache.scala 525:49]
  wire [22:0] a_mask; // @[DCache.scala 529:29]
  wire [2:0] _T_1412; // @[Misc.scala 201:34]
  wire [3:0] _T_1414; // @[OneHot.scala 65:12]
  wire [2:0] _T_1416; // @[Misc.scala 201:81]
  wire  _T_1417; // @[Misc.scala 205:21]
  wire  _T_1422; // @[Misc.scala 214:38]
  wire  _T_1423; // @[Misc.scala 214:29]
  wire  _T_1425; // @[Misc.scala 214:38]
  wire  _T_1426; // @[Misc.scala 214:29]
  wire  _T_1430; // @[Misc.scala 213:27]
  wire  _T_1431; // @[Misc.scala 214:38]
  wire  _T_1432; // @[Misc.scala 214:29]
  wire  _T_1433; // @[Misc.scala 213:27]
  wire  _T_1434; // @[Misc.scala 214:38]
  wire  _T_1435; // @[Misc.scala 214:29]
  wire  _T_1436; // @[Misc.scala 213:27]
  wire  _T_1437; // @[Misc.scala 214:38]
  wire  _T_1438; // @[Misc.scala 214:29]
  wire  _T_1439; // @[Misc.scala 213:27]
  wire  _T_1440; // @[Misc.scala 214:38]
  wire  _T_1441; // @[Misc.scala 214:29]
  wire  _T_1445; // @[Misc.scala 213:27]
  wire  _T_1446; // @[Misc.scala 214:38]
  wire  _T_1447; // @[Misc.scala 214:29]
  wire  _T_1448; // @[Misc.scala 213:27]
  wire  _T_1449; // @[Misc.scala 214:38]
  wire  _T_1450; // @[Misc.scala 214:29]
  wire  _T_1451; // @[Misc.scala 213:27]
  wire  _T_1452; // @[Misc.scala 214:38]
  wire  _T_1453; // @[Misc.scala 214:29]
  wire  _T_1454; // @[Misc.scala 213:27]
  wire  _T_1455; // @[Misc.scala 214:38]
  wire  _T_1456; // @[Misc.scala 214:29]
  wire  _T_1457; // @[Misc.scala 213:27]
  wire  _T_1458; // @[Misc.scala 214:38]
  wire  _T_1459; // @[Misc.scala 214:29]
  wire  _T_1460; // @[Misc.scala 213:27]
  wire  _T_1461; // @[Misc.scala 214:38]
  wire  _T_1462; // @[Misc.scala 214:29]
  wire  _T_1463; // @[Misc.scala 213:27]
  wire  _T_1464; // @[Misc.scala 214:38]
  wire  _T_1465; // @[Misc.scala 214:29]
  wire  _T_1466; // @[Misc.scala 213:27]
  wire  _T_1467; // @[Misc.scala 214:38]
  wire  _T_1468; // @[Misc.scala 214:29]
  wire [7:0] get_mask; // @[Cat.scala 29:58]
  wire  _T_2577; // @[Mux.scala 80:60]
  wire [2:0] _T_2578_opcode; // @[Mux.scala 80:57]
  wire [3:0] _T_1696_size; // @[Edges.scala 515:17 Edges.scala 518:15]
  wire [3:0] _T_2578_size; // @[Mux.scala 80:57]
  wire  _T_2578_source; // @[Mux.scala 80:57]
  wire [31:0] _T_2578_address; // @[Mux.scala 80:57]
  wire [7:0] _T_2578_mask; // @[Mux.scala 80:57]
  wire [63:0] _T_2578_data; // @[Mux.scala 80:57]
  wire  _T_2579; // @[Mux.scala 80:60]
  wire [2:0] _T_2580_opcode; // @[Mux.scala 80:57]
  wire [2:0] _T_2580_param; // @[Mux.scala 80:57]
  wire [3:0] _T_2580_size; // @[Mux.scala 80:57]
  wire  _T_2580_source; // @[Mux.scala 80:57]
  wire [31:0] _T_2580_address; // @[Mux.scala 80:57]
  wire [7:0] _T_2580_mask; // @[Mux.scala 80:57]
  wire [63:0] _T_2580_data; // @[Mux.scala 80:57]
  wire  _T_2581; // @[Mux.scala 80:60]
  wire [2:0] _T_2582_opcode; // @[Mux.scala 80:57]
  wire [2:0] _T_2582_param; // @[Mux.scala 80:57]
  wire [3:0] _T_2582_size; // @[Mux.scala 80:57]
  wire  _T_2582_source; // @[Mux.scala 80:57]
  wire [31:0] _T_2582_address; // @[Mux.scala 80:57]
  wire [7:0] _T_2582_mask; // @[Mux.scala 80:57]
  wire [63:0] _T_2582_data; // @[Mux.scala 80:57]
  wire  _T_2583; // @[Mux.scala 80:60]
  wire [2:0] _T_2584_opcode; // @[Mux.scala 80:57]
  wire [2:0] _T_2584_param; // @[Mux.scala 80:57]
  wire [3:0] _T_2584_size; // @[Mux.scala 80:57]
  wire  _T_2584_source; // @[Mux.scala 80:57]
  wire [31:0] _T_2584_address; // @[Mux.scala 80:57]
  wire [7:0] _T_2584_mask; // @[Mux.scala 80:57]
  wire [63:0] _T_2584_data; // @[Mux.scala 80:57]
  wire  _T_2585; // @[Mux.scala 80:60]
  wire [2:0] _T_2586_opcode; // @[Mux.scala 80:57]
  wire [2:0] _T_2586_param; // @[Mux.scala 80:57]
  wire [3:0] _T_2586_size; // @[Mux.scala 80:57]
  wire  _T_2586_source; // @[Mux.scala 80:57]
  wire [31:0] _T_2586_address; // @[Mux.scala 80:57]
  wire [7:0] _T_2586_mask; // @[Mux.scala 80:57]
  wire [63:0] _T_2586_data; // @[Mux.scala 80:57]
  wire  _T_2587; // @[Mux.scala 80:60]
  wire [2:0] _T_2588_opcode; // @[Mux.scala 80:57]
  wire [2:0] _T_2588_param; // @[Mux.scala 80:57]
  wire [3:0] _T_2588_size; // @[Mux.scala 80:57]
  wire  _T_2588_source; // @[Mux.scala 80:57]
  wire [31:0] _T_2588_address; // @[Mux.scala 80:57]
  wire [7:0] _T_2588_mask; // @[Mux.scala 80:57]
  wire [63:0] _T_2588_data; // @[Mux.scala 80:57]
  wire  _T_2589; // @[Mux.scala 80:60]
  wire [2:0] _T_2590_opcode; // @[Mux.scala 80:57]
  wire [2:0] _T_2590_param; // @[Mux.scala 80:57]
  wire [3:0] _T_2590_size; // @[Mux.scala 80:57]
  wire  _T_2590_source; // @[Mux.scala 80:57]
  wire [31:0] _T_2590_address; // @[Mux.scala 80:57]
  wire [7:0] _T_2590_mask; // @[Mux.scala 80:57]
  wire [63:0] _T_2590_data; // @[Mux.scala 80:57]
  wire  _T_2591; // @[Mux.scala 80:60]
  wire [2:0] _T_2592_opcode; // @[Mux.scala 80:57]
  wire [2:0] _T_2592_param; // @[Mux.scala 80:57]
  wire [3:0] _T_2592_size; // @[Mux.scala 80:57]
  wire  _T_2592_source; // @[Mux.scala 80:57]
  wire [31:0] _T_2592_address; // @[Mux.scala 80:57]
  wire [7:0] _T_2592_mask; // @[Mux.scala 80:57]
  wire [63:0] _T_2592_data; // @[Mux.scala 80:57]
  wire  _T_2593; // @[Mux.scala 80:60]
  wire [2:0] atomics_opcode; // @[Mux.scala 80:57]
  wire [2:0] atomics_param; // @[Mux.scala 80:57]
  wire [3:0] atomics_size; // @[Mux.scala 80:57]
  wire  atomics_source; // @[Mux.scala 80:57]
  wire [31:0] atomics_address; // @[Mux.scala 80:57]
  wire [7:0] atomics_mask; // @[Mux.scala 80:57]
  wire [63:0] atomics_data; // @[Mux.scala 80:57]
  wire  _T_2596; // @[DCache.scala 551:27]
  wire  _T_2600; // @[DCache.scala 551:48]
  wire  tl_out_a_valid; // @[DCache.scala 550:67]
  wire [2:0] _T_2693_opcode; // @[DCache.scala 555:8]
  wire [2:0] _T_2693_param; // @[DCache.scala 555:8]
  wire [3:0] _T_2693_size; // @[DCache.scala 555:8]
  wire  _T_2693_source; // @[DCache.scala 555:8]
  wire [31:0] _T_2693_address; // @[DCache.scala 555:8]
  wire [7:0] _T_2693_mask; // @[DCache.scala 555:8]
  wire [63:0] _T_2693_data; // @[DCache.scala 555:8]
  wire [2:0] _T_2694_opcode; // @[DCache.scala 554:8]
  wire [2:0] _T_2694_param; // @[DCache.scala 554:8]
  wire [3:0] _T_2694_size; // @[DCache.scala 554:8]
  wire  _T_2694_source; // @[DCache.scala 554:8]
  wire [31:0] _T_2694_address; // @[DCache.scala 554:8]
  wire [7:0] putpartial_mask; // @[Edges.scala 485:17 Edges.scala 491:15]
  wire [7:0] _T_2694_mask; // @[DCache.scala 554:8]
  wire [63:0] _T_2694_data; // @[DCache.scala 554:8]
  wire [2:0] _T_2695_opcode; // @[DCache.scala 553:8]
  wire [2:0] _T_2695_param; // @[DCache.scala 553:8]
  wire [3:0] _T_2695_size; // @[DCache.scala 553:8]
  wire  _T_2695_source; // @[DCache.scala 553:8]
  wire [31:0] _T_2695_address; // @[DCache.scala 553:8]
  wire [7:0] _T_2695_mask; // @[DCache.scala 553:8]
  wire [63:0] _T_2695_data; // @[DCache.scala 553:8]
  wire [2:0] _T_2625_param; // @[Edges.scala 347:17 Edges.scala 349:15]
  wire [1:0] _T_2698; // @[OneHot.scala 65:12]
  wire  a_sel; // @[DCache.scala 574:66]
  wire  _T_2700; // @[Decoupled.scala 40:37]
  wire  _GEN_143; // @[DCache.scala 578:18]
  wire [26:0] _T_2707; // @[package.scala 212:77]
  wire [8:0] _T_2710; // @[Edges.scala 221:59]
  wire [8:0] _T_2712; // @[Edges.scala 222:14]
  wire [8:0] _T_2715; // @[Edges.scala 231:28]
  wire  _T_2716; // @[Edges.scala 233:25]
  wire  _T_2717; // @[Edges.scala 233:47]
  wire  d_last; // @[Edges.scala 233:37]
  wire  d_done; // @[Edges.scala 234:22]
  wire [8:0] _T_2719; // @[Edges.scala 235:25]
  wire [11:0] d_address_inc; // @[Edges.scala 270:29]
  wire  grantIsVoluntary; // @[DCache.scala 608:32]
  wire [2:0] _T_2749; // @[DCache.scala 612:97]
  wire [1:0] _T_2758; // @[OneHot.scala 65:12]
  wire  uncachedRespIdxOH; // @[DCache.scala 615:90]
  wire  _T_2763; // @[DCache.scala 620:13]
  wire  _T_2766; // @[DCache.scala 629:17]
  wire  _T_2768; // @[DCache.scala 630:17]
  wire [31:0] dontCareBits; // @[DCache.scala 644:55]
  wire [31:0] _GEN_347; // @[DCache.scala 645:26]
  wire [31:0] _T_2773; // @[DCache.scala 645:26]
  wire  _T_2775; // @[DCache.scala 651:13]
  wire  _GEN_195; // @[DCache.scala 650:36]
  wire  _GEN_204; // @[DCache.scala 627:35]
  wire  _GEN_208; // @[DCache.scala 618:26]
  wire  _GEN_217; // @[DCache.scala 618:26]
  wire  _GEN_230; // @[DCache.scala 617:26]
  wire  _T_2777; // @[DCache.scala 657:36]
  wire  _T_2778; // @[DCache.scala 657:47]
  wire  _T_2779; // @[DCache.scala 657:64]
  wire  tl_out__e_valid; // @[DCache.scala 665:51]
  wire  _T_2781; // @[Decoupled.scala 40:37]
  wire  _T_2783; // @[DCache.scala 659:47]
  wire  _T_2784; // @[DCache.scala 659:58]
  wire  _T_2785; // @[DCache.scala 659:26]
  wire  _T_2787; // @[DCache.scala 659:9]
  wire  _T_2789; // @[DCache.scala 664:44]
  wire  _T_2790; // @[DCache.scala 664:61]
  wire [39:0] _T_2794; // @[DCache.scala 671:57]
  wire [39:0] _GEN_348; // @[DCache.scala 671:67]
  wire [39:0] _T_2795; // @[DCache.scala 671:67]
  wire  _T_2798; // @[DCache.scala 684:43]
  wire [3:0] _T_2857; // @[Cat.scala 29:58]
  wire  _T_2866; // @[Mux.scala 80:60]
  wire [1:0] _T_2867; // @[Mux.scala 80:57]
  wire  _T_2868; // @[Mux.scala 80:60]
  wire [1:0] _T_2869; // @[Mux.scala 80:57]
  wire  _T_2870; // @[Mux.scala 80:60]
  wire [1:0] _T_2871; // @[Mux.scala 80:57]
  wire  _T_2872; // @[Mux.scala 80:60]
  wire [1:0] _T_2873; // @[Mux.scala 80:57]
  wire  _GEN_233; // @[DCache.scala 698:29]
  wire  _GEN_234; // @[DCache.scala 698:29]
  wire  _GEN_235; // @[DCache.scala 698:29]
  wire  _T_2888; // @[DCache.scala 712:79]
  wire  _T_2889; // @[DCache.scala 712:44]
  wire [39:0] _T_2897; // @[Cat.scala 29:58]
  wire [8:0] _T_2908; // @[Edges.scala 231:28]
  wire [8:0] c_count; // @[Edges.scala 235:25]
  reg  s1_release_data_valid; // @[DCache.scala 723:34]
  reg [31:0] _RAND_92;
  wire  releaseRejected; // @[DCache.scala 725:44]
  wire [9:0] _T_2919; // @[Cat.scala 29:58]
  wire [1:0] _T_2920; // @[Cat.scala 29:58]
  wire [1:0] _GEN_349; // @[DCache.scala 726:101]
  wire [1:0] _T_2922; // @[DCache.scala 726:101]
  wire [1:0] _T_2923; // @[DCache.scala 726:52]
  wire [9:0] _GEN_350; // @[DCache.scala 726:47]
  wire [9:0] releaseDataBeat; // @[DCache.scala 726:47]
  wire  _T_2928; // @[DCache.scala 739:34]
  wire  _T_2929; // @[DCache.scala 739:52]
  wire  _T_2931; // @[DCache.scala 739:13]
  wire  discard_line; // @[DCache.scala 740:46]
  wire  _T_2938; // @[DCache.scala 741:44]
  wire [2:0] _T_2939; // @[DCache.scala 741:27]
  wire [25:0] _T_2941; // @[Cat.scala 29:58]
  wire [31:0] res_2_address; // @[DCache.scala 742:96]
  wire [2:0] _GEN_243; // @[DCache.scala 738:25]
  wire [2:0] _T_2944; // @[DCache.scala 753:29]
  wire [2:0] _T_2946; // @[DCache.scala 757:29]
  wire [2:0] _GEN_254; // @[DCache.scala 750:45]
  wire [2:0] _GEN_260; // @[DCache.scala 750:45]
  wire [2:0] _GEN_262; // @[DCache.scala 748:36]
  wire [2:0] _GEN_265; // @[DCache.scala 748:36]
  wire [2:0] _GEN_272; // @[DCache.scala 746:28]
  wire [2:0] _GEN_275; // @[DCache.scala 746:28]
  wire [2:0] _GEN_283; // @[DCache.scala 744:21]
  wire [2:0] _GEN_286; // @[DCache.scala 744:21]
  wire  _T_2947; // @[DCache.scala 761:25]
  wire [39:0] _T_2950; // @[Cat.scala 29:58]
  wire [2:0] _GEN_293; // @[DCache.scala 765:37]
  wire  _GEN_294; // @[DCache.scala 765:37]
  wire [2:0] _GEN_298; // @[DCache.scala 761:44]
  wire [2:0] _GEN_300; // @[DCache.scala 772:26]
  wire [2:0] _GEN_302; // @[DCache.scala 770:47]
  wire [2:0] _GEN_306; // @[DCache.scala 774:48]
  wire [2:0] _GEN_315; // @[DCache.scala 779:48]
  wire  _T_2978; // @[DCache.scala 792:29]
  wire  _GEN_323; // @[DCache.scala 792:41]
  wire [1:0] newCoh_state; // @[DCache.scala 783:81]
  wire  _T_2980; // @[DCache.scala 803:60]
  wire [11:0] _T_2983; // @[DCache.scala 806:55]
  wire [5:0] _T_2985; // @[DCache.scala 806:117]
  wire [11:0] _GEN_352; // @[DCache.scala 806:72]
  wire  _T_2990; // @[package.scala 15:47]
  wire  _T_2999; // @[Decoupled.scala 40:37]
  wire  _T_3006; // @[DCache.scala 829:57]
  wire  _T_3007; // @[DCache.scala 829:94]
  wire  _T_3009; // @[DCache.scala 829:115]
  wire  _T_3012; // @[DCache.scala 831:40]
  reg  _T_3014; // @[DCache.scala 832:32]
  reg [31:0] _RAND_93;
  reg  doUncachedResp; // @[DCache.scala 847:27]
  reg [31:0] _RAND_94;
  wire  _T_3027; // @[DCache.scala 851:11]
  wire [31:0] _T_3035; // @[AMOALU.scala 39:24]
  wire  _T_3038; // @[AMOALU.scala 42:26]
  wire  _T_3041; // @[AMOALU.scala 42:76]
  wire [31:0] _T_3043; // @[Bitwise.scala 72:12]
  wire [31:0] _T_3045; // @[AMOALU.scala 42:20]
  wire [63:0] _T_3046; // @[Cat.scala 29:58]
  wire [15:0] _T_3050; // @[AMOALU.scala 39:24]
  wire  _T_3053; // @[AMOALU.scala 42:26]
  wire  _T_3056; // @[AMOALU.scala 42:76]
  wire [47:0] _T_3058; // @[Bitwise.scala 72:12]
  wire [47:0] _T_3060; // @[AMOALU.scala 42:20]
  wire [63:0] _T_3061; // @[Cat.scala 29:58]
  wire [7:0] _T_3065; // @[AMOALU.scala 39:24]
  wire [7:0] _T_3067; // @[AMOALU.scala 41:23]
  wire  _T_3068; // @[AMOALU.scala 42:26]
  wire  _T_3069; // @[AMOALU.scala 42:38]
  wire  _T_3071; // @[AMOALU.scala 42:76]
  wire [55:0] _T_3073; // @[Bitwise.scala 72:12]
  wire [55:0] _T_3075; // @[AMOALU.scala 42:20]
  wire [63:0] _T_3076; // @[Cat.scala 29:58]
  wire [63:0] _GEN_353; // @[DCache.scala 873:41]
  reg  resetting; // @[DCache.scala 906:26]
  reg [31:0] _RAND_95;
  reg  _T_3097; // @[DCache.scala 908:18]
  reg [31:0] _RAND_96;
  wire  _GEN_341; // @[DCache.scala 908:27]
  reg [7:0] flushCounter; // @[DCache.scala 909:25]
  reg [31:0] _RAND_97;
  wire [8:0] flushCounterNext; // @[DCache.scala 910:39]
  wire  flushDone; // @[DCache.scala 911:57]
  wire  _T_3103; // @[Decoupled.scala 40:37]
  wire  _T_3105; // @[DCache.scala 915:45]
  wire  _T_3107; // @[DCache.scala 915:64]
  wire  _T_3109; // @[DCache.scala 915:95]
  wire [11:0] _T_3116; // @[DCache.scala 919:98]
  wire [8:0] _GEN_343; // @[DCache.scala 952:20]
  reg [8:0] _T_3178; // @[Edges.scala 230:27]
  reg [31:0] _RAND_98;
  wire [8:0] _T_3180; // @[Edges.scala 231:28]
  wire  _T_3181; // @[Edges.scala 232:25]
  wire  _T_3182; // @[Edges.scala 233:25]
  wire  _T_3184; // @[Edges.scala 233:37]
  wire  _GEN_356; // @[DCache.scala 620:13]
  wire  _GEN_359; // @[DCache.scala 630:17]
  wire  _GEN_360; // @[DCache.scala 630:17]
  wire  _GEN_361; // @[DCache.scala 630:17]
  wire  _GEN_369; // @[DCache.scala 651:13]
  wire  _GEN_370; // @[DCache.scala 651:13]
  reg [19:0] DCache_state; // @[Register tracking DCache state]
  reg [31:0] _RAND_99;
  reg  DCache_cov [0:1048575]; // @[Coverage map for DCache]
  reg [31:0] _RAND_100;
  wire  DCache_cov_read_data; // @[Coverage map for DCache]
  wire [19:0] DCache_cov_read_addr; // @[Coverage map for DCache]
  wire  DCache_cov_write_data; // @[Coverage map for DCache]
  wire [19:0] DCache_cov_write_addr; // @[Coverage map for DCache]
  wire  DCache_cov_write_mask; // @[Coverage map for DCache]
  wire  DCache_cov_write_en; // @[Coverage map for DCache]
  reg [29:0] DCache_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_101;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire [9:0] pstore1_held_shl;
  wire [19:0] pstore1_held_pad;
  wire [5:0] pstore2_valid_shl;
  wire [19:0] pstore2_valid_pad;
  wire [2:0] s2_valid_shl;
  wire [19:0] s2_valid_pad;
  wire [17:0] release_state_shl;
  wire [19:0] release_state_pad;
  wire [7:0] s2_probe_shl;
  wire [19:0] s2_probe_pad;
  wire  s2_flush_valid_pre_tag_ecc_shl;
  wire [19:0] s2_flush_valid_pre_tag_ecc_pad;
  wire [10:0] _T_679_state_shl;
  wire [19:0] _T_679_state_pad;
  wire [1:0] uncachedInFlight_0_shl;
  wire [19:0] uncachedInFlight_0_pad;
  wire [14:0] s2_release_data_valid_shl;
  wire [19:0] s2_release_data_valid_pad;
  wire [7:0] probe_bits_param_shl;
  wire [19:0] probe_bits_param_pad;
  wire [14:0] s2_pma_cacheable_shl;
  wire [19:0] s2_pma_cacheable_pad;
  wire [13:0] s2_hit_state_state_shl;
  wire [19:0] s2_hit_state_state_pad;
  wire [1:0] s2_req_size_shl;
  wire [19:0] s2_req_size_pad;
  wire  s1_did_read_shl;
  wire [19:0] s1_did_read_pad;
  wire [11:0] grantInProgress_shl;
  wire [19:0] grantInProgress_pad;
  wire [11:0] _T_1016_shl;
  wire [19:0] _T_1016_pad;
  wire [12:0] s2_not_nacked_in_s1_shl;
  wire [19:0] s2_not_nacked_in_s1_pad;
  wire [19:0] blockUncachedGrant_shl;
  wire [19:0] blockUncachedGrant_pad;
  wire [16:0] _T_672_shl;
  wire [19:0] _T_672_pad;
  wire [6:0] s2_hit_way_shl;
  wire [19:0] s2_hit_way_pad;
  wire [19:0] cached_grant_wait_shl;
  wire [19:0] cached_grant_wait_pad;
  wire [11:0] s2_req_signed_shl;
  wire [19:0] s2_req_signed_pad;
  wire [16:0] release_ack_wait_shl;
  wire [19:0] release_ack_wait_pad;
  wire [3:0] s2_probe_state_state_shl;
  wire [19:0] s2_probe_state_state_pad;
  wire [2:0] s1_probe_shl;
  wire [19:0] s1_probe_pad;
  wire [1:0] s1_valid_shl;
  wire [19:0] s1_valid_pad;
  wire [6:0] s1_req_size_shl;
  wire [19:0] s1_req_size_pad;
  wire [15:0] pstore1_rmw_shl;
  wire [19:0] pstore1_rmw_pad;
  wire [11:0] s1_flush_valid_shl;
  wire [19:0] s1_flush_valid_pad;
  wire  resetting_shl;
  wire [19:0] resetting_pad;
  wire [15:0] s2_probe_way_shl;
  wire [19:0] s2_probe_way_pad;
  wire [9:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [2:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [7:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [15:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [5:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [19:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [19:0] DCache_xor15;
  wire [19:0] DCache_xor16;
  wire [19:0] DCache_xor7;
  wire [19:0] DCache_xor17;
  wire [19:0] DCache_xor38;
  wire [19:0] DCache_xor18;
  wire [19:0] DCache_xor8;
  wire [19:0] DCache_xor3;
  wire [19:0] DCache_xor19;
  wire [19:0] DCache_xor20;
  wire [19:0] DCache_xor9;
  wire [19:0] DCache_xor21;
  wire [19:0] DCache_xor46;
  wire [19:0] DCache_xor22;
  wire [19:0] DCache_xor10;
  wire [19:0] DCache_xor4;
  wire [19:0] DCache_xor1;
  wire [19:0] DCache_xor23;
  wire [19:0] DCache_xor24;
  wire [19:0] DCache_xor11;
  wire [19:0] DCache_xor25;
  wire [19:0] DCache_xor54;
  wire [19:0] DCache_xor26;
  wire [19:0] DCache_xor12;
  wire [19:0] DCache_xor5;
  wire [19:0] DCache_xor27;
  wire [19:0] DCache_xor58;
  wire [19:0] DCache_xor28;
  wire [19:0] DCache_xor13;
  wire [19:0] DCache_xor29;
  wire [19:0] DCache_xor62;
  wire [19:0] DCache_xor30;
  wire [19:0] DCache_xor14;
  wire [19:0] DCache_xor6;
  wire [19:0] DCache_xor2;
  wire [19:0] DCache_xor0;
  wire [29:0] amoalu_sum;
  wire [29:0] MaxPeriodFibonacciLFSR_sum;
  wire [29:0] pma_checker_sum;
  wire [29:0] metaArb_sum;
  wire [29:0] dataArb_sum;
  wire [29:0] tlb_sum;
  wire [29:0] data_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  stopEn4;
  wire  stopEn5;
  wire  stopEn6;
  wire  stopEn7;
  wire  stopEn8;
  wire  stopEn9;
  wire  MaxPeriodFibonacciLFSR_metaAssert_wire;
  wire  dataArb_metaAssert_wire;
  wire  metaArb_metaAssert_wire;
  wire  tlb_metaAssert_wire;
  wire  pma_checker_metaAssert_wire;
  wire  data_metaAssert_wire;
  wire  amoalu_metaAssert_wire;
  wire  DCache_or7;
  wire  DCache_or8;
  wire  DCache_or3;
  wire  DCache_or9;
  wire  DCache_or10;
  wire  DCache_or4;
  wire  DCache_or1;
  wire  DCache_or11;
  wire  DCache_or12;
  wire  DCache_or5;
  wire  DCache_or13;
  wire  DCache_or30;
  wire  DCache_or14;
  wire  DCache_or6;
  wire  DCache_or2;
  wire  DCache_or0;
  TLB tlb ( // @[DCache.scala 115:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vaddr(tlb_io_req_bits_vaddr),
    .io_req_bits_passthrough(tlb_io_req_bits_passthrough),
    .io_req_bits_size(tlb_io_req_bits_size),
    .io_req_bits_cmd(tlb_io_req_bits_cmd),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_paddr(tlb_io_resp_paddr),
    .io_resp_pf_ld(tlb_io_resp_pf_ld),
    .io_resp_pf_st(tlb_io_resp_pf_st),
    .io_resp_ae_ld(tlb_io_resp_ae_ld),
    .io_resp_ae_st(tlb_io_resp_ae_st),
    .io_resp_ma_ld(tlb_io_resp_ma_ld),
    .io_resp_ma_st(tlb_io_resp_ma_st),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_sfence_valid(tlb_io_sfence_valid),
    .io_sfence_bits_rs1(tlb_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(tlb_io_sfence_bits_rs2),
    .io_sfence_bits_addr(tlb_io_sfence_bits_addr),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_bits_addr(tlb_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(tlb_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(tlb_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(tlb_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(tlb_io_ptw_ptbr_mode),
    .io_ptw_status_debug(tlb_io_ptw_status_debug),
    .io_ptw_status_dprv(tlb_io_ptw_status_dprv),
    .io_ptw_status_mxr(tlb_io_ptw_status_mxr),
    .io_ptw_status_sum(tlb_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(tlb_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(tlb_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(tlb_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(tlb_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(tlb_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(tlb_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(tlb_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(tlb_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(tlb_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(tlb_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(tlb_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(tlb_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(tlb_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(tlb_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(tlb_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(tlb_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(tlb_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(tlb_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(tlb_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(tlb_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(tlb_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(tlb_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(tlb_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(tlb_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(tlb_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(tlb_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(tlb_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(tlb_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(tlb_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(tlb_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(tlb_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(tlb_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(tlb_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(tlb_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(tlb_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(tlb_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(tlb_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(tlb_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(tlb_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(tlb_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(tlb_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(tlb_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(tlb_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(tlb_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(tlb_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(tlb_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(tlb_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(tlb_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(tlb_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(tlb_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(tlb_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(tlb_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(tlb_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(tlb_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(tlb_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(tlb_io_ptw_pmp_7_mask),
    .io_covSum(tlb_io_covSum),
    .metaAssert(tlb_metaAssert),
    .metaReset(tlb_metaReset)
  );
  TLB pma_checker ( // @[DCache.scala 116:27]
    .clock(pma_checker_clock),
    .reset(pma_checker_reset),
    .io_req_ready(pma_checker_io_req_ready),
    .io_req_valid(pma_checker_io_req_valid),
    .io_req_bits_vaddr(pma_checker_io_req_bits_vaddr),
    .io_req_bits_passthrough(pma_checker_io_req_bits_passthrough),
    .io_req_bits_size(pma_checker_io_req_bits_size),
    .io_req_bits_cmd(pma_checker_io_req_bits_cmd),
    .io_resp_miss(pma_checker_io_resp_miss),
    .io_resp_paddr(pma_checker_io_resp_paddr),
    .io_resp_pf_ld(pma_checker_io_resp_pf_ld),
    .io_resp_pf_st(pma_checker_io_resp_pf_st),
    .io_resp_ae_ld(pma_checker_io_resp_ae_ld),
    .io_resp_ae_st(pma_checker_io_resp_ae_st),
    .io_resp_ma_ld(pma_checker_io_resp_ma_ld),
    .io_resp_ma_st(pma_checker_io_resp_ma_st),
    .io_resp_cacheable(pma_checker_io_resp_cacheable),
    .io_sfence_valid(pma_checker_io_sfence_valid),
    .io_sfence_bits_rs1(pma_checker_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(pma_checker_io_sfence_bits_rs2),
    .io_sfence_bits_addr(pma_checker_io_sfence_bits_addr),
    .io_ptw_req_ready(pma_checker_io_ptw_req_ready),
    .io_ptw_req_valid(pma_checker_io_ptw_req_valid),
    .io_ptw_req_bits_bits_addr(pma_checker_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(pma_checker_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(pma_checker_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(pma_checker_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(pma_checker_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(pma_checker_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(pma_checker_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(pma_checker_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(pma_checker_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(pma_checker_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(pma_checker_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(pma_checker_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(pma_checker_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(pma_checker_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(pma_checker_io_ptw_ptbr_mode),
    .io_ptw_status_debug(pma_checker_io_ptw_status_debug),
    .io_ptw_status_dprv(pma_checker_io_ptw_status_dprv),
    .io_ptw_status_mxr(pma_checker_io_ptw_status_mxr),
    .io_ptw_status_sum(pma_checker_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(pma_checker_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(pma_checker_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(pma_checker_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(pma_checker_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(pma_checker_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(pma_checker_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(pma_checker_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(pma_checker_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(pma_checker_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(pma_checker_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(pma_checker_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(pma_checker_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(pma_checker_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(pma_checker_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(pma_checker_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(pma_checker_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(pma_checker_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(pma_checker_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(pma_checker_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(pma_checker_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(pma_checker_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(pma_checker_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(pma_checker_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(pma_checker_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(pma_checker_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(pma_checker_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(pma_checker_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(pma_checker_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(pma_checker_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(pma_checker_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(pma_checker_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(pma_checker_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(pma_checker_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(pma_checker_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(pma_checker_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(pma_checker_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(pma_checker_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(pma_checker_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(pma_checker_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(pma_checker_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(pma_checker_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(pma_checker_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(pma_checker_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(pma_checker_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(pma_checker_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(pma_checker_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(pma_checker_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(pma_checker_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(pma_checker_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(pma_checker_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(pma_checker_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(pma_checker_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(pma_checker_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(pma_checker_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(pma_checker_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(pma_checker_io_ptw_pmp_7_mask),
    .io_covSum(pma_checker_io_covSum),
    .metaAssert(pma_checker_metaAssert),
    .metaReset(pma_checker_metaReset)
  );
  MaxPeriodFibonacciLFSR MaxPeriodFibonacciLFSR ( // @[PRNG.scala 82:22]
    .clock(MaxPeriodFibonacciLFSR_clock),
    .reset(MaxPeriodFibonacciLFSR_reset),
    .io_increment(MaxPeriodFibonacciLFSR_io_increment),
    .io_out_0(MaxPeriodFibonacciLFSR_io_out_0),
    .io_out_1(MaxPeriodFibonacciLFSR_io_out_1),
    .io_out_2(MaxPeriodFibonacciLFSR_io_out_2),
    .io_out_3(MaxPeriodFibonacciLFSR_io_out_3),
    .io_out_4(MaxPeriodFibonacciLFSR_io_out_4),
    .io_out_5(MaxPeriodFibonacciLFSR_io_out_5),
    .io_out_6(MaxPeriodFibonacciLFSR_io_out_6),
    .io_out_7(MaxPeriodFibonacciLFSR_io_out_7),
    .io_out_8(MaxPeriodFibonacciLFSR_io_out_8),
    .io_out_9(MaxPeriodFibonacciLFSR_io_out_9),
    .io_out_10(MaxPeriodFibonacciLFSR_io_out_10),
    .io_out_11(MaxPeriodFibonacciLFSR_io_out_11),
    .io_out_12(MaxPeriodFibonacciLFSR_io_out_12),
    .io_out_13(MaxPeriodFibonacciLFSR_io_out_13),
    .io_out_14(MaxPeriodFibonacciLFSR_io_out_14),
    .io_out_15(MaxPeriodFibonacciLFSR_io_out_15),
    .io_covSum(MaxPeriodFibonacciLFSR_io_covSum),
    .metaAssert(MaxPeriodFibonacciLFSR_metaAssert),
    .metaReset(MaxPeriodFibonacciLFSR_metaReset)
  );
  DCacheModuleImpl_Anon_1 metaArb ( // @[DCache.scala 120:23]
    .io_in_0_valid(metaArb_io_in_0_valid),
    .io_in_0_bits_addr(metaArb_io_in_0_bits_addr),
    .io_in_0_bits_idx(metaArb_io_in_0_bits_idx),
    .io_in_0_bits_data(metaArb_io_in_0_bits_data),
    .io_in_1_valid(metaArb_io_in_1_valid),
    .io_in_1_bits_addr(metaArb_io_in_1_bits_addr),
    .io_in_1_bits_idx(metaArb_io_in_1_bits_idx),
    .io_in_1_bits_data(metaArb_io_in_1_bits_data),
    .io_in_2_valid(metaArb_io_in_2_valid),
    .io_in_2_bits_addr(metaArb_io_in_2_bits_addr),
    .io_in_2_bits_idx(metaArb_io_in_2_bits_idx),
    .io_in_2_bits_way_en(metaArb_io_in_2_bits_way_en),
    .io_in_2_bits_data(metaArb_io_in_2_bits_data),
    .io_in_3_valid(metaArb_io_in_3_valid),
    .io_in_3_bits_addr(metaArb_io_in_3_bits_addr),
    .io_in_3_bits_idx(metaArb_io_in_3_bits_idx),
    .io_in_3_bits_way_en(metaArb_io_in_3_bits_way_en),
    .io_in_3_bits_data(metaArb_io_in_3_bits_data),
    .io_in_4_ready(metaArb_io_in_4_ready),
    .io_in_4_valid(metaArb_io_in_4_valid),
    .io_in_4_bits_addr(metaArb_io_in_4_bits_addr),
    .io_in_4_bits_idx(metaArb_io_in_4_bits_idx),
    .io_in_4_bits_way_en(metaArb_io_in_4_bits_way_en),
    .io_in_4_bits_data(metaArb_io_in_4_bits_data),
    .io_in_5_ready(metaArb_io_in_5_ready),
    .io_in_5_valid(metaArb_io_in_5_valid),
    .io_in_5_bits_addr(metaArb_io_in_5_bits_addr),
    .io_in_5_bits_idx(metaArb_io_in_5_bits_idx),
    .io_in_6_ready(metaArb_io_in_6_ready),
    .io_in_6_valid(metaArb_io_in_6_valid),
    .io_in_6_bits_addr(metaArb_io_in_6_bits_addr),
    .io_in_6_bits_idx(metaArb_io_in_6_bits_idx),
    .io_in_6_bits_way_en(metaArb_io_in_6_bits_way_en),
    .io_in_6_bits_data(metaArb_io_in_6_bits_data),
    .io_in_7_ready(metaArb_io_in_7_ready),
    .io_in_7_valid(metaArb_io_in_7_valid),
    .io_in_7_bits_addr(metaArb_io_in_7_bits_addr),
    .io_in_7_bits_idx(metaArb_io_in_7_bits_idx),
    .io_in_7_bits_way_en(metaArb_io_in_7_bits_way_en),
    .io_in_7_bits_data(metaArb_io_in_7_bits_data),
    .io_out_valid(metaArb_io_out_valid),
    .io_out_bits_write(metaArb_io_out_bits_write),
    .io_out_bits_addr(metaArb_io_out_bits_addr),
    .io_out_bits_idx(metaArb_io_out_bits_idx),
    .io_out_bits_way_en(metaArb_io_out_bits_way_en),
    .io_out_bits_data(metaArb_io_out_bits_data),
    .io_covSum(metaArb_io_covSum),
    .metaAssert(metaArb_metaAssert)
  );
  DCacheDataArray data ( // @[DCache.scala 130:20]
    .clock(data_clock),
    .io_req_valid(data_io_req_valid),
    .io_req_bits_addr(data_io_req_bits_addr),
    .io_req_bits_write(data_io_req_bits_write),
    .io_req_bits_wdata(data_io_req_bits_wdata),
    .io_req_bits_eccMask(data_io_req_bits_eccMask),
    .io_req_bits_way_en(data_io_req_bits_way_en),
    .io_resp_0(data_io_resp_0),
    .io_resp_1(data_io_resp_1),
    .io_resp_2(data_io_resp_2),
    .io_resp_3(data_io_resp_3),
    .io_covSum(data_io_covSum),
    .metaAssert(data_metaAssert),
    .metaReset(data_metaReset)
  );
  DCacheModuleImpl_Anon_2 dataArb ( // @[DCache.scala 131:23]
    .io_in_0_valid(dataArb_io_in_0_valid),
    .io_in_0_bits_addr(dataArb_io_in_0_bits_addr),
    .io_in_0_bits_write(dataArb_io_in_0_bits_write),
    .io_in_0_bits_wdata(dataArb_io_in_0_bits_wdata),
    .io_in_0_bits_eccMask(dataArb_io_in_0_bits_eccMask),
    .io_in_0_bits_way_en(dataArb_io_in_0_bits_way_en),
    .io_in_1_ready(dataArb_io_in_1_ready),
    .io_in_1_valid(dataArb_io_in_1_valid),
    .io_in_1_bits_addr(dataArb_io_in_1_bits_addr),
    .io_in_1_bits_write(dataArb_io_in_1_bits_write),
    .io_in_1_bits_wdata(dataArb_io_in_1_bits_wdata),
    .io_in_1_bits_eccMask(dataArb_io_in_1_bits_eccMask),
    .io_in_1_bits_way_en(dataArb_io_in_1_bits_way_en),
    .io_in_2_ready(dataArb_io_in_2_ready),
    .io_in_2_valid(dataArb_io_in_2_valid),
    .io_in_2_bits_addr(dataArb_io_in_2_bits_addr),
    .io_in_2_bits_wdata(dataArb_io_in_2_bits_wdata),
    .io_in_2_bits_eccMask(dataArb_io_in_2_bits_eccMask),
    .io_in_3_ready(dataArb_io_in_3_ready),
    .io_in_3_valid(dataArb_io_in_3_valid),
    .io_in_3_bits_addr(dataArb_io_in_3_bits_addr),
    .io_in_3_bits_wdata(dataArb_io_in_3_bits_wdata),
    .io_in_3_bits_eccMask(dataArb_io_in_3_bits_eccMask),
    .io_out_valid(dataArb_io_out_valid),
    .io_out_bits_addr(dataArb_io_out_bits_addr),
    .io_out_bits_write(dataArb_io_out_bits_write),
    .io_out_bits_wdata(dataArb_io_out_bits_wdata),
    .io_out_bits_eccMask(dataArb_io_out_bits_eccMask),
    .io_out_bits_way_en(dataArb_io_out_bits_way_en),
    .io_covSum(dataArb_io_covSum),
    .metaAssert(dataArb_metaAssert)
  );
  AMOALU amoalu ( // @[DCache.scala 881:26]
    .io_mask(amoalu_io_mask),
    .io_cmd(amoalu_io_cmd),
    .io_lhs(amoalu_io_lhs),
    .io_rhs(amoalu_io_rhs),
    .io_out(amoalu_io_out),
    .io_covSum(amoalu_io_covSum),
    .metaAssert(amoalu_metaAssert)
  );
  assign tag_array_0_s1_meta_addr = tag_array_0_s1_meta_addr_pipe_0;
  assign tag_array_0_s1_meta_data = tag_array_0[tag_array_0_s1_meta_addr]; // @[DescribedSRAM.scala 23:26]
  assign tag_array_0__T_260_data = metaArb_io_out_bits_data;
  assign tag_array_0__T_260_addr = metaArb_io_out_bits_idx;
  assign tag_array_0__T_260_mask = metaArb_io_out_bits_way_en[0];
  assign tag_array_0__T_260_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign tag_array_1_s1_meta_addr = tag_array_1_s1_meta_addr_pipe_0;
  assign tag_array_1_s1_meta_data = tag_array_1[tag_array_1_s1_meta_addr]; // @[DescribedSRAM.scala 23:26]
  assign tag_array_1__T_260_data = metaArb_io_out_bits_data;
  assign tag_array_1__T_260_addr = metaArb_io_out_bits_idx;
  assign tag_array_1__T_260_mask = metaArb_io_out_bits_way_en[1];
  assign tag_array_1__T_260_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign tag_array_2_s1_meta_addr = tag_array_2_s1_meta_addr_pipe_0;
  assign tag_array_2_s1_meta_data = tag_array_2[tag_array_2_s1_meta_addr]; // @[DescribedSRAM.scala 23:26]
  assign tag_array_2__T_260_data = metaArb_io_out_bits_data;
  assign tag_array_2__T_260_addr = metaArb_io_out_bits_idx;
  assign tag_array_2__T_260_mask = metaArb_io_out_bits_way_en[2];
  assign tag_array_2__T_260_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign tag_array_3_s1_meta_addr = tag_array_3_s1_meta_addr_pipe_0;
  assign tag_array_3_s1_meta_data = tag_array_3[tag_array_3_s1_meta_addr]; // @[DescribedSRAM.scala 23:26]
  assign tag_array_3__T_260_data = metaArb_io_out_bits_data;
  assign tag_array_3__T_260_addr = metaArb_io_out_bits_idx;
  assign tag_array_3__T_260_mask = metaArb_io_out_bits_way_en[3];
  assign tag_array_3__T_260_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign _T_7 = {MaxPeriodFibonacciLFSR_io_out_7,MaxPeriodFibonacciLFSR_io_out_6,MaxPeriodFibonacciLFSR_io_out_5,MaxPeriodFibonacciLFSR_io_out_4,MaxPeriodFibonacciLFSR_io_out_3,MaxPeriodFibonacciLFSR_io_out_2,MaxPeriodFibonacciLFSR_io_out_1,MaxPeriodFibonacciLFSR_io_out_0}; // @[PRNG.scala 86:17]
  assign _T_15 = {MaxPeriodFibonacciLFSR_io_out_15,MaxPeriodFibonacciLFSR_io_out_14,MaxPeriodFibonacciLFSR_io_out_13,MaxPeriodFibonacciLFSR_io_out_12,MaxPeriodFibonacciLFSR_io_out_11,MaxPeriodFibonacciLFSR_io_out_10,MaxPeriodFibonacciLFSR_io_out_9,MaxPeriodFibonacciLFSR_io_out_8,_T_7}; // @[PRNG.scala 86:17]
  assign _T_16 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  assign _T_2882 = blockProbeAfterGrantCount > 3'h0; // @[DCache.scala 709:65]
  assign lrscValid = lrscCount > 7'h3; // @[DCache.scala 424:29]
  assign block_probe_for_core_progress = _T_2882 | lrscValid; // @[DCache.scala 709:69]
  assign _T_381 = s1_probe | s2_probe; // @[DCache.scala 286:34]
  assign _T_382 = release_state != 3'h0; // @[DCache.scala 286:63]
  assign releaseInFlight = _T_381 | _T_382; // @[DCache.scala 286:46]
  assign _T_2883 = auto_out_b_bits_address ^ release_ack_addr; // @[DCache.scala 710:88]
  assign _T_2885 = _T_2883[11:6] == 6'h0; // @[DCache.scala 710:124]
  assign block_probe_for_pending_release_ack = release_ack_wait & _T_2885; // @[DCache.scala 710:62]
  assign _T_2886 = releaseInFlight | block_probe_for_pending_release_ack; // @[DCache.scala 711:50]
  assign block_probe_for_ordering = _T_2886 | grantInProgress; // @[DCache.scala 711:89]
  assign _T_2890 = block_probe_for_core_progress | block_probe_for_ordering; // @[DCache.scala 713:79]
  assign _T_2891 = _T_2890 | s1_valid; // @[DCache.scala 713:107]
  assign _T_2892 = _T_2891 | s2_valid; // @[DCache.scala 713:119]
  assign tl_out__b_ready = metaArb_io_in_6_ready & ~_T_2892; // @[DCache.scala 713:44]
  assign _T_17 = tl_out__b_ready & auto_out_b_valid; // @[Decoupled.scala 40:37]
  assign s1_valid_masked = s1_valid & ~io_cpu_s1_kill; // @[DCache.scala 163:34]
  assign s2_meta_error = |4'h0; // @[DCache.scala 314:83]
  assign _T_680 = {probe_bits_param,s2_probe_state_state}; // @[Cat.scala 29:58]
  assign _T_737 = 4'h3 == _T_680; // @[Misc.scala 55:20]
  assign _T_733 = 4'h2 == _T_680; // @[Misc.scala 55:20]
  assign _T_729 = 4'h1 == _T_680; // @[Misc.scala 55:20]
  assign _T_725 = 4'h0 == _T_680; // @[Misc.scala 55:20]
  assign _T_721 = 4'h7 == _T_680; // @[Misc.scala 55:20]
  assign _T_717 = 4'h6 == _T_680; // @[Misc.scala 55:20]
  assign _T_713 = 4'h5 == _T_680; // @[Misc.scala 55:20]
  assign _T_709 = 4'h4 == _T_680; // @[Misc.scala 55:20]
  assign _T_705 = 4'hb == _T_680; // @[Misc.scala 55:20]
  assign _T_701 = 4'ha == _T_680; // @[Misc.scala 55:20]
  assign _T_697 = 4'h9 == _T_680; // @[Misc.scala 55:20]
  assign _T_693 = 4'h8 == _T_680; // @[Misc.scala 55:20]
  assign _T_710 = _T_709 ? 1'h0 : _T_705; // @[Misc.scala 37:9]
  assign _T_714 = _T_713 ? 1'h0 : _T_710; // @[Misc.scala 37:9]
  assign _T_718 = _T_717 ? 1'h0 : _T_714; // @[Misc.scala 37:9]
  assign _T_722 = _T_721 | _T_718; // @[Misc.scala 37:9]
  assign _T_726 = _T_725 ? 1'h0 : _T_722; // @[Misc.scala 37:9]
  assign _T_730 = _T_729 ? 1'h0 : _T_726; // @[Misc.scala 37:9]
  assign _T_734 = _T_733 ? 1'h0 : _T_730; // @[Misc.scala 37:9]
  assign s2_prb_ack_data = _T_737 | _T_734; // @[Misc.scala 37:9]
  assign _T_2943 = s2_probe_state_state > 2'h0; // @[Metadata.scala 50:45]
  assign _T_2909 = _T_2906 == 9'h1; // @[Edges.scala 233:25]
  assign _T_2954 = release_state == 3'h1; // @[package.scala 15:47]
  assign _T_2955 = release_state == 3'h6; // @[package.scala 15:47]
  assign _T_2956 = _T_2954 | _T_2955; // @[package.scala 64:59]
  assign _T_2953 = release_state == 3'h2; // @[DCache.scala 779:25]
  assign _T_2952 = release_state == 3'h3; // @[DCache.scala 774:25]
  assign _GEN_314 = _T_2953 ? 3'h5 : 3'h4; // @[DCache.scala 779:48]
  assign tl_out__c_bits_opcode = _T_2956 ? 3'h7 : _GEN_314; // @[DCache.scala 783:81]
  assign tl_out__c_bits_size = _T_2956 ? 4'h6 : probe_bits_size; // @[DCache.scala 783:81]
  assign _T_2900 = 27'hfff << tl_out__c_bits_size; // @[package.scala 212:77]
  assign _T_2903 = ~_T_2900[11:3]; // @[Edges.scala 221:59]
  assign _T_2905 = tl_out__c_bits_opcode[0] ? _T_2903 : 9'h0; // @[Edges.scala 222:14]
  assign _T_2910 = _T_2905 == 9'h0; // @[Edges.scala 233:47]
  assign c_last = _T_2909 | _T_2910; // @[Edges.scala 233:37]
  assign _T_2951 = release_state == 3'h5; // @[DCache.scala 770:25]
  assign c_first = _T_2906 == 9'h0; // @[Edges.scala 232:25]
  assign _T_2925 = c_first & release_ack_wait; // @[DCache.scala 732:56]
  assign _T_2927 = s2_release_data_valid & ~_T_2925; // @[DCache.scala 732:43]
  assign _GEN_263 = s2_prb_ack_data ? _T_2927 : 1'h1; // @[DCache.scala 748:36]
  assign _GEN_273 = s2_meta_error ? _T_2927 : _GEN_263; // @[DCache.scala 746:28]
  assign _GEN_284 = s2_probe ? _GEN_273 : _T_2927; // @[DCache.scala 744:21]
  assign _GEN_301 = _T_2951 | _GEN_284; // @[DCache.scala 770:47]
  assign tl_out__c_valid = _T_2952 | _GEN_301; // @[DCache.scala 774:48]
  assign _T_2898 = auto_out_c_ready & tl_out__c_valid; // @[Decoupled.scala 40:37]
  assign releaseDone = c_last & _T_2898; // @[Edges.scala 234:22]
  assign _GEN_261 = _T_2943 | ~releaseDone; // @[DCache.scala 750:45]
  assign _GEN_271 = s2_prb_ack_data | _GEN_261; // @[DCache.scala 748:36]
  assign probeNack = s2_meta_error | _GEN_271; // @[DCache.scala 746:28]
  assign _T_30 = s1_req_cmd == 5'h0; // @[Consts.scala 82:31]
  assign _T_31 = s1_req_cmd == 5'h6; // @[Consts.scala 82:48]
  assign _T_32 = _T_30 | _T_31; // @[Consts.scala 82:41]
  assign _T_33 = s1_req_cmd == 5'h7; // @[Consts.scala 82:65]
  assign _T_34 = _T_32 | _T_33; // @[Consts.scala 82:58]
  assign _T_35 = s1_req_cmd == 5'h4; // @[package.scala 15:47]
  assign _T_36 = s1_req_cmd == 5'h9; // @[package.scala 15:47]
  assign _T_39 = _T_35 | _T_36; // @[package.scala 64:59]
  assign _T_37 = s1_req_cmd == 5'ha; // @[package.scala 15:47]
  assign _T_40 = _T_39 | _T_37; // @[package.scala 64:59]
  assign _T_38 = s1_req_cmd == 5'hb; // @[package.scala 15:47]
  assign _T_41 = _T_40 | _T_38; // @[package.scala 64:59]
  assign _T_42 = s1_req_cmd == 5'h8; // @[package.scala 15:47]
  assign _T_43 = s1_req_cmd == 5'hc; // @[package.scala 15:47]
  assign _T_47 = _T_42 | _T_43; // @[package.scala 64:59]
  assign _T_44 = s1_req_cmd == 5'hd; // @[package.scala 15:47]
  assign _T_48 = _T_47 | _T_44; // @[package.scala 64:59]
  assign _T_45 = s1_req_cmd == 5'he; // @[package.scala 15:47]
  assign _T_49 = _T_48 | _T_45; // @[package.scala 64:59]
  assign _T_46 = s1_req_cmd == 5'hf; // @[package.scala 15:47]
  assign _T_50 = _T_49 | _T_46; // @[package.scala 64:59]
  assign _T_51 = _T_41 | _T_50; // @[Consts.scala 80:44]
  assign s1_read = _T_34 | _T_51; // @[Consts.scala 82:75]
  assign _T_418 = s2_req_cmd == 5'h1; // @[Consts.scala 83:32]
  assign _T_419 = s2_req_cmd == 5'h11; // @[Consts.scala 83:49]
  assign _T_420 = _T_418 | _T_419; // @[Consts.scala 83:42]
  assign _T_421 = s2_req_cmd == 5'h7; // @[Consts.scala 83:66]
  assign _T_422 = _T_420 | _T_421; // @[Consts.scala 83:59]
  assign _T_423 = s2_req_cmd == 5'h4; // @[package.scala 15:47]
  assign _T_424 = s2_req_cmd == 5'h9; // @[package.scala 15:47]
  assign _T_427 = _T_423 | _T_424; // @[package.scala 64:59]
  assign _T_425 = s2_req_cmd == 5'ha; // @[package.scala 15:47]
  assign _T_428 = _T_427 | _T_425; // @[package.scala 64:59]
  assign _T_426 = s2_req_cmd == 5'hb; // @[package.scala 15:47]
  assign _T_429 = _T_428 | _T_426; // @[package.scala 64:59]
  assign _T_430 = s2_req_cmd == 5'h8; // @[package.scala 15:47]
  assign _T_431 = s2_req_cmd == 5'hc; // @[package.scala 15:47]
  assign _T_435 = _T_430 | _T_431; // @[package.scala 64:59]
  assign _T_432 = s2_req_cmd == 5'hd; // @[package.scala 15:47]
  assign _T_436 = _T_435 | _T_432; // @[package.scala 64:59]
  assign _T_433 = s2_req_cmd == 5'he; // @[package.scala 15:47]
  assign _T_437 = _T_436 | _T_433; // @[package.scala 64:59]
  assign _T_434 = s2_req_cmd == 5'hf; // @[package.scala 15:47]
  assign _T_438 = _T_437 | _T_434; // @[package.scala 64:59]
  assign _T_439 = _T_429 | _T_438; // @[Consts.scala 80:44]
  assign s2_write = _T_422 | _T_439; // @[Consts.scala 83:76]
  assign _T_1017 = s2_valid & s2_write; // @[DCache.scala 456:39]
  assign pstore1_valid_likely = _T_1017 | pstore1_held; // @[DCache.scala 456:51]
  assign _T_1178 = pstore1_addr[11:3] == s1_req_addr[11:3]; // @[DCache.scala 508:31]
  assign _T_52 = s1_req_cmd == 5'h1; // @[Consts.scala 83:32]
  assign _T_53 = s1_req_cmd == 5'h11; // @[Consts.scala 83:49]
  assign _T_54 = _T_52 | _T_53; // @[Consts.scala 83:42]
  assign _T_56 = _T_54 | _T_33; // @[Consts.scala 83:59]
  assign s1_write = _T_56 | _T_51; // @[Consts.scala 83:76]
  assign _T_1194 = |pstore1_mask[7]; // @[DCache.scala 1076:66]
  assign _T_1193 = |pstore1_mask[6]; // @[DCache.scala 1076:66]
  assign _T_1192 = |pstore1_mask[5]; // @[DCache.scala 1076:66]
  assign _T_1191 = |pstore1_mask[4]; // @[DCache.scala 1076:66]
  assign _T_1190 = |pstore1_mask[3]; // @[DCache.scala 1076:66]
  assign _T_1189 = |pstore1_mask[2]; // @[DCache.scala 1076:66]
  assign _T_1188 = |pstore1_mask[1]; // @[DCache.scala 1076:66]
  assign _T_1187 = |pstore1_mask[0]; // @[DCache.scala 1076:66]
  assign _T_1201 = {_T_1194,_T_1193,_T_1192,_T_1191,_T_1190,_T_1189,_T_1188,_T_1187}; // @[Cat.scala 29:58]
  assign _T_1216 = {_T_1201[7],_T_1201[6],_T_1201[5],_T_1201[4],_T_1201[3],_T_1201[2],_T_1201[1],_T_1201[0]}; // @[Cat.scala 29:58]
  assign _T_340 = s1_req_size >= 2'h1; // @[AMOALU.scala 17:57]
  assign _T_342 = s1_req_addr[0] | _T_340; // @[AMOALU.scala 17:46]
  assign _T_344 = s1_req_addr[0] ? 1'h0 : 1'h1; // @[AMOALU.scala 18:22]
  assign _T_345 = {_T_342,_T_344}; // @[Cat.scala 29:58]
  assign _T_347 = s1_req_addr[1] ? _T_345 : 2'h0; // @[AMOALU.scala 17:22]
  assign _T_348 = s1_req_size >= 2'h2; // @[AMOALU.scala 17:57]
  assign _T_349 = _T_348 ? 2'h3 : 2'h0; // @[AMOALU.scala 17:51]
  assign _T_350 = _T_347 | _T_349; // @[AMOALU.scala 17:46]
  assign _T_352 = s1_req_addr[1] ? 2'h0 : _T_345; // @[AMOALU.scala 18:22]
  assign _T_353 = {_T_350,_T_352}; // @[Cat.scala 29:58]
  assign _T_355 = s1_req_addr[2] ? _T_353 : 4'h0; // @[AMOALU.scala 17:22]
  assign _T_356 = s1_req_size >= 2'h3; // @[AMOALU.scala 17:57]
  assign _T_357 = _T_356 ? 4'hf : 4'h0; // @[AMOALU.scala 17:51]
  assign _T_358 = _T_355 | _T_357; // @[AMOALU.scala 17:46]
  assign _T_360 = s1_req_addr[2] ? 4'h0 : _T_353; // @[AMOALU.scala 18:22]
  assign s1_mask_xwr = {_T_358,_T_360}; // @[Cat.scala 29:58]
  assign _T_1232 = |s1_mask_xwr[7]; // @[DCache.scala 1076:66]
  assign _T_1231 = |s1_mask_xwr[6]; // @[DCache.scala 1076:66]
  assign _T_1230 = |s1_mask_xwr[5]; // @[DCache.scala 1076:66]
  assign _T_1229 = |s1_mask_xwr[4]; // @[DCache.scala 1076:66]
  assign _T_1228 = |s1_mask_xwr[3]; // @[DCache.scala 1076:66]
  assign _T_1227 = |s1_mask_xwr[2]; // @[DCache.scala 1076:66]
  assign _T_1226 = |s1_mask_xwr[1]; // @[DCache.scala 1076:66]
  assign _T_1225 = |s1_mask_xwr[0]; // @[DCache.scala 1076:66]
  assign _T_1239 = {_T_1232,_T_1231,_T_1230,_T_1229,_T_1228,_T_1227,_T_1226,_T_1225}; // @[Cat.scala 29:58]
  assign _T_1254 = {_T_1239[7],_T_1239[6],_T_1239[5],_T_1239[4],_T_1239[3],_T_1239[2],_T_1239[1],_T_1239[0]}; // @[Cat.scala 29:58]
  assign _T_1255 = _T_1216 & _T_1254; // @[DCache.scala 509:38]
  assign _T_1256 = |_T_1255; // @[DCache.scala 509:66]
  assign _T_1257 = pstore1_mask & s1_mask_xwr; // @[DCache.scala 509:77]
  assign _T_1258 = |_T_1257; // @[DCache.scala 509:92]
  assign _T_1259 = s1_write ? _T_1256 : _T_1258; // @[DCache.scala 509:8]
  assign _T_1260 = _T_1178 & _T_1259; // @[DCache.scala 508:68]
  assign _T_1261 = pstore1_valid_likely & _T_1260; // @[DCache.scala 511:27]
  assign _T_1264 = pstore2_addr[11:3] == s1_req_addr[11:3]; // @[DCache.scala 508:31]
  assign _T_1280 = |mask[7]; // @[DCache.scala 1076:66]
  assign _T_1279 = |mask[6]; // @[DCache.scala 1076:66]
  assign _T_1278 = |mask[5]; // @[DCache.scala 1076:66]
  assign _T_1277 = |mask[4]; // @[DCache.scala 1076:66]
  assign _T_1276 = |mask[3]; // @[DCache.scala 1076:66]
  assign _T_1275 = |mask[2]; // @[DCache.scala 1076:66]
  assign _T_1274 = |mask[1]; // @[DCache.scala 1076:66]
  assign _T_1273 = |mask[0]; // @[DCache.scala 1076:66]
  assign _T_1287 = {_T_1280,_T_1279,_T_1278,_T_1277,_T_1276,_T_1275,_T_1274,_T_1273}; // @[Cat.scala 29:58]
  assign _T_1302 = {_T_1287[7],_T_1287[6],_T_1287[5],_T_1287[4],_T_1287[3],_T_1287[2],_T_1287[1],_T_1287[0]}; // @[Cat.scala 29:58]
  assign _T_1341 = _T_1302 & _T_1254; // @[DCache.scala 509:38]
  assign _T_1342 = |_T_1341; // @[DCache.scala 509:66]
  assign _T_1343 = mask & s1_mask_xwr; // @[DCache.scala 509:77]
  assign _T_1344 = |_T_1343; // @[DCache.scala 509:92]
  assign _T_1345 = s1_write ? _T_1342 : _T_1344; // @[DCache.scala 509:8]
  assign _T_1346 = _T_1264 & _T_1345; // @[DCache.scala 508:68]
  assign _T_1347 = pstore2_valid & _T_1346; // @[DCache.scala 512:21]
  assign s1_hazard = _T_1261 | _T_1347; // @[DCache.scala 511:69]
  assign s1_raw_hazard = s1_read & s1_hazard; // @[DCache.scala 513:31]
  assign _T_1348 = s1_valid & s1_raw_hazard; // @[DCache.scala 518:18]
  assign _T_378 = {io_cpu_s2_xcpt_ma_ld,io_cpu_s2_xcpt_ma_st,io_cpu_s2_xcpt_pf_ld,io_cpu_s2_xcpt_pf_st,io_cpu_s2_xcpt_ae_ld,io_cpu_s2_xcpt_ae_st}; // @[DCache.scala 284:54]
  assign _T_379 = |_T_378; // @[DCache.scala 284:61]
  assign s2_valid_no_xcpt = s2_valid & ~_T_379; // @[DCache.scala 284:35]
  assign s2_valid_masked = s2_valid_no_xcpt & s2_not_nacked_in_s1; // @[DCache.scala 289:42]
  assign _T_644 = s2_valid_masked & ~s2_meta_error; // @[DCache.scala 349:71]
  assign _T_539 = s2_req_cmd == 5'h3; // @[Consts.scala 84:54]
  assign _T_540 = s2_write | _T_539; // @[Consts.scala 84:47]
  assign _T_541 = s2_req_cmd == 5'h6; // @[Consts.scala 84:71]
  assign _T_542 = _T_540 | _T_541; // @[Consts.scala 84:64]
  assign _T_544 = {s2_write,_T_542,s2_hit_state_state}; // @[Cat.scala 29:58]
  assign _T_602 = 4'h3 == _T_544; // @[Misc.scala 48:20]
  assign _T_599 = 4'h2 == _T_544; // @[Misc.scala 48:20]
  assign _T_596 = 4'h1 == _T_544; // @[Misc.scala 48:20]
  assign _T_593 = 4'h7 == _T_544; // @[Misc.scala 48:20]
  assign _T_590 = 4'h6 == _T_544; // @[Misc.scala 48:20]
  assign _T_587 = 4'hf == _T_544; // @[Misc.scala 48:20]
  assign _T_584 = 4'he == _T_544; // @[Misc.scala 48:20]
  assign _T_581 = 4'h0 == _T_544; // @[Misc.scala 48:20]
  assign _T_578 = 4'h5 == _T_544; // @[Misc.scala 48:20]
  assign _T_575 = 4'h4 == _T_544; // @[Misc.scala 48:20]
  assign _T_572 = 4'hd == _T_544; // @[Misc.scala 48:20]
  assign _T_569 = 4'hc == _T_544; // @[Misc.scala 48:20]
  assign _T_588 = _T_587 | _T_584; // @[Misc.scala 34:9]
  assign _T_591 = _T_590 | _T_588; // @[Misc.scala 34:9]
  assign _T_594 = _T_593 | _T_591; // @[Misc.scala 34:9]
  assign _T_597 = _T_596 | _T_594; // @[Misc.scala 34:9]
  assign _T_600 = _T_599 | _T_597; // @[Misc.scala 34:9]
  assign s2_hit = _T_602 | _T_600; // @[Misc.scala 34:9]
  assign s2_valid_hit_maybe_flush_pre_data_ecc_and_waw = _T_644 & s2_hit; // @[DCache.scala 349:89]
  assign _T_396 = s2_req_cmd == 5'h0; // @[Consts.scala 82:31]
  assign _T_398 = _T_396 | _T_541; // @[Consts.scala 82:41]
  assign _T_400 = _T_398 | _T_421; // @[Consts.scala 82:58]
  assign s2_read = _T_400 | _T_439; // @[Consts.scala 82:75]
  assign s2_readwrite = s2_read | s2_write; // @[DCache.scala 306:30]
  assign s2_valid_hit_pre_data_ecc_and_waw = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_readwrite; // @[DCache.scala 370:89]
  assign _T_571 = _T_569 ? 2'h1 : 2'h0; // @[Misc.scala 34:36]
  assign _T_574 = _T_572 ? 2'h2 : _T_571; // @[Misc.scala 34:36]
  assign _T_577 = _T_575 ? 2'h1 : _T_574; // @[Misc.scala 34:36]
  assign _T_580 = _T_578 ? 2'h2 : _T_577; // @[Misc.scala 34:36]
  assign _T_583 = _T_581 ? 2'h0 : _T_580; // @[Misc.scala 34:36]
  assign _T_586 = _T_584 ? 2'h3 : _T_583; // @[Misc.scala 34:36]
  assign _T_589 = _T_587 ? 2'h3 : _T_586; // @[Misc.scala 34:36]
  assign _T_592 = _T_590 ? 2'h2 : _T_589; // @[Misc.scala 34:36]
  assign _T_595 = _T_593 ? 2'h3 : _T_592; // @[Misc.scala 34:36]
  assign _T_598 = _T_596 ? 2'h1 : _T_595; // @[Misc.scala 34:36]
  assign _T_601 = _T_599 ? 2'h2 : _T_598; // @[Misc.scala 34:36]
  assign s2_grow_param = _T_602 ? 2'h3 : _T_601; // @[Misc.scala 34:36]
  assign _T_804 = s2_hit_state_state == s2_grow_param; // @[Metadata.scala 46:46]
  assign s2_update_meta = ~_T_804; // @[Metadata.scala 47:40]
  assign _T_823 = s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta; // @[DCache.scala 397:62]
  assign _T_824 = io_cpu_s2_nack | _T_823; // @[DCache.scala 397:24]
  assign s1_readwrite = s1_read | s1_write; // @[DCache.scala 185:30]
  assign _T_74 = s1_req_cmd == 5'h5; // @[DCache.scala 187:34]
  assign s1_flush_line = _T_74 & s1_req_size[0]; // @[DCache.scala 187:50]
  assign _T_227 = s1_readwrite | s1_flush_line; // @[DCache.scala 229:38]
  assign _T_228 = s1_req_cmd == 5'h17; // @[DCache.scala 229:69]
  assign s1_cmd_uses_tlb = _T_227 | _T_228; // @[DCache.scala 229:55]
  assign _T_242 = s1_valid & s1_cmd_uses_tlb; // @[DCache.scala 235:39]
  assign _T_243 = _T_242 & tlb_io_resp_miss; // @[DCache.scala 235:58]
  assign _GEN_118 = _T_824 | _T_243; // @[DCache.scala 397:82]
  assign _GEN_142 = _T_1348 | _GEN_118; // @[DCache.scala 518:36]
  assign _GEN_282 = probeNack | _GEN_142; // @[DCache.scala 759:24]
  assign s1_nack = s2_probe ? _GEN_282 : _GEN_142; // @[DCache.scala 744:21]
  assign s1_valid_not_nacked = s1_valid & ~s1_nack; // @[DCache.scala 164:38]
  assign s0_clk_en = metaArb_io_out_valid & ~metaArb_io_out_bits_write; // @[DCache.scala 167:40]
  assign s0_req_addr = {metaArb_io_out_bits_addr[39:6],io_cpu_req_bits_addr[5:0]}; // @[Cat.scala 29:58]
  assign s0_req_phys = ~metaArb_io_in_7_ready | io_cpu_req_bits_phys; // @[DCache.scala 171:34]
  assign s1_sfence = s1_req_cmd == 5'h14; // @[DCache.scala 186:30]
  assign inWriteback = _T_2954 | _T_2953; // @[package.scala 64:59]
  assign _T_78 = release_state == 3'h0; // @[DCache.scala 203:38]
  assign _T_80 = _T_78 & ~cached_grant_wait; // @[DCache.scala 203:51]
  assign _T_82 = _T_80 & ~s1_nack; // @[DCache.scala 203:73]
  assign _T_84 = io_cpu_req_bits_cmd == 5'h0; // @[Consts.scala 82:31]
  assign _T_85 = io_cpu_req_bits_cmd == 5'h6; // @[Consts.scala 82:48]
  assign _T_86 = _T_84 | _T_85; // @[Consts.scala 82:41]
  assign _T_87 = io_cpu_req_bits_cmd == 5'h7; // @[Consts.scala 82:65]
  assign _T_88 = _T_86 | _T_87; // @[Consts.scala 82:58]
  assign _T_89 = io_cpu_req_bits_cmd == 5'h4; // @[package.scala 15:47]
  assign _T_90 = io_cpu_req_bits_cmd == 5'h9; // @[package.scala 15:47]
  assign _T_91 = io_cpu_req_bits_cmd == 5'ha; // @[package.scala 15:47]
  assign _T_92 = io_cpu_req_bits_cmd == 5'hb; // @[package.scala 15:47]
  assign _T_93 = _T_89 | _T_90; // @[package.scala 64:59]
  assign _T_94 = _T_93 | _T_91; // @[package.scala 64:59]
  assign _T_95 = _T_94 | _T_92; // @[package.scala 64:59]
  assign _T_96 = io_cpu_req_bits_cmd == 5'h8; // @[package.scala 15:47]
  assign _T_97 = io_cpu_req_bits_cmd == 5'hc; // @[package.scala 15:47]
  assign _T_98 = io_cpu_req_bits_cmd == 5'hd; // @[package.scala 15:47]
  assign _T_99 = io_cpu_req_bits_cmd == 5'he; // @[package.scala 15:47]
  assign _T_100 = io_cpu_req_bits_cmd == 5'hf; // @[package.scala 15:47]
  assign _T_101 = _T_96 | _T_97; // @[package.scala 64:59]
  assign _T_102 = _T_101 | _T_98; // @[package.scala 64:59]
  assign _T_103 = _T_102 | _T_99; // @[package.scala 64:59]
  assign _T_104 = _T_103 | _T_100; // @[package.scala 64:59]
  assign _T_105 = _T_95 | _T_104; // @[Consts.scala 80:44]
  assign s0_read = _T_88 | _T_105; // @[Consts.scala 82:75]
  assign _T_106 = io_cpu_req_bits_cmd == 5'h1; // @[package.scala 15:47]
  assign _T_107 = io_cpu_req_bits_cmd == 5'h3; // @[package.scala 15:47]
  assign _T_108 = _T_106 | _T_107; // @[package.scala 64:59]
  assign res = ~_T_108; // @[DCache.scala 1080:15]
  assign _T_135 = io_cpu_req_bits_cmd == 5'h11; // @[Consts.scala 83:49]
  assign _T_136 = _T_106 | _T_135; // @[Consts.scala 83:42]
  assign _T_138 = _T_136 | _T_87; // @[Consts.scala 83:59]
  assign _T_156 = _T_138 | _T_105; // @[Consts.scala 83:76]
  assign _T_160 = _T_156 & _T_135; // @[DCache.scala 1086:23]
  assign _T_161 = s0_read | _T_160; // @[DCache.scala 1085:21]
  assign _T_163 = ~_T_161 | res; // @[DCache.scala 1081:28]
  assign _T_165 = _T_163 | reset; // @[DCache.scala 1081:11]
  assign _T_167 = io_cpu_req_valid & res; // @[DCache.scala 212:46]
  assign _T_171 = ~dataArb_io_in_3_ready & s0_read; // @[DCache.scala 218:33]
  assign _GEN_28 = _T_171 ? 1'h0 : _T_82; // @[DCache.scala 218:45]
  assign _T_223 = io_cpu_req_valid & _T_161; // @[DCache.scala 219:75]
  assign _T_224 = dataArb_io_in_3_ready & _T_223; // @[DCache.scala 219:54]
  assign _GEN_30 = metaArb_io_in_7_ready ? _GEN_28 : 1'h0; // @[DCache.scala 226:34]
  assign _T_237 = ~tlb_io_req_ready & ~tlb_io_ptw_resp_valid; // @[DCache.scala 234:27]
  assign _T_239 = _T_237 & ~io_cpu_req_bits_phys; // @[DCache.scala 234:53]
  assign _GEN_31 = _T_239 ? 1'h0 : _GEN_30; // @[DCache.scala 234:79]
  assign s1_paddr = {tlb_io_resp_paddr[31:12],s1_req_addr[11:0]}; // @[Cat.scala 29:58]
  assign s1_victim_way = _T_15[1:0]; // @[package.scala 143:13]
  assign _T_266 = tag_array_0_s1_meta_data;
  assign s1_meta_uncorrected_0_tag = _T_266[19:0]; // @[DCache.scala 267:80]
  assign s1_meta_uncorrected_0_coh_state = _T_266[21:20]; // @[DCache.scala 267:80]
  assign _T_269 = tag_array_1_s1_meta_data;
  assign s1_meta_uncorrected_1_tag = _T_269[19:0]; // @[DCache.scala 267:80]
  assign s1_meta_uncorrected_1_coh_state = _T_269[21:20]; // @[DCache.scala 267:80]
  assign _T_272 = tag_array_2_s1_meta_data;
  assign s1_meta_uncorrected_2_tag = _T_272[19:0]; // @[DCache.scala 267:80]
  assign s1_meta_uncorrected_2_coh_state = _T_272[21:20]; // @[DCache.scala 267:80]
  assign _T_275 = tag_array_3_s1_meta_data;
  assign s1_meta_uncorrected_3_tag = _T_275[19:0]; // @[DCache.scala 267:80]
  assign s1_meta_uncorrected_3_coh_state = _T_275[21:20]; // @[DCache.scala 267:80]
  assign s1_tag = s1_paddr[31:12]; // @[DCache.scala 268:29]
  assign _T_278 = s1_meta_uncorrected_0_coh_state > 2'h0; // @[Metadata.scala 50:45]
  assign _T_279 = s1_meta_uncorrected_0_tag == s1_tag; // @[DCache.scala 269:83]
  assign _T_280 = _T_278 & _T_279; // @[DCache.scala 269:74]
  assign _T_281 = s1_meta_uncorrected_1_coh_state > 2'h0; // @[Metadata.scala 50:45]
  assign _T_282 = s1_meta_uncorrected_1_tag == s1_tag; // @[DCache.scala 269:83]
  assign _T_283 = _T_281 & _T_282; // @[DCache.scala 269:74]
  assign _T_284 = s1_meta_uncorrected_2_coh_state > 2'h0; // @[Metadata.scala 50:45]
  assign _T_285 = s1_meta_uncorrected_2_tag == s1_tag; // @[DCache.scala 269:83]
  assign _T_286 = _T_284 & _T_285; // @[DCache.scala 269:74]
  assign _T_287 = s1_meta_uncorrected_3_coh_state > 2'h0; // @[Metadata.scala 50:45]
  assign _T_288 = s1_meta_uncorrected_3_tag == s1_tag; // @[DCache.scala 269:83]
  assign _T_289 = _T_287 & _T_288; // @[DCache.scala 269:74]
  assign s1_meta_hit_way = {_T_289,_T_286,_T_283,_T_280}; // @[Cat.scala 29:58]
  assign _T_295 = _T_279 & ~s1_flush_valid; // @[DCache.scala 271:59]
  assign _T_296 = _T_295 ? s1_meta_uncorrected_0_coh_state : 2'h0; // @[DCache.scala 271:41]
  assign _T_299 = _T_282 & ~s1_flush_valid; // @[DCache.scala 271:59]
  assign _T_300 = _T_299 ? s1_meta_uncorrected_1_coh_state : 2'h0; // @[DCache.scala 271:41]
  assign _T_303 = _T_285 & ~s1_flush_valid; // @[DCache.scala 271:59]
  assign _T_304 = _T_303 ? s1_meta_uncorrected_2_coh_state : 2'h0; // @[DCache.scala 271:41]
  assign _T_307 = _T_288 & ~s1_flush_valid; // @[DCache.scala 271:59]
  assign _T_308 = _T_307 ? s1_meta_uncorrected_3_coh_state : 2'h0; // @[DCache.scala 271:41]
  assign _T_309 = _T_296 | _T_300; // @[DCache.scala 272:19]
  assign _T_310 = _T_309 | _T_304; // @[DCache.scala 272:19]
  assign s1_meta_hit_state_state = _T_310 | _T_308; // @[DCache.scala 272:19]
  assign _T_316 = s1_victim_way == 2'h1; // @[package.scala 32:86]
  assign _T_318 = s1_victim_way == 2'h2; // @[package.scala 32:86]
  assign _T_320 = s1_victim_way == 2'h3; // @[package.scala 32:86]
  assign s2_hit_valid = s2_hit_state_state > 2'h0; // @[Metadata.scala 50:45]
  assign _T_673 = 4'h1 << _T_672; // @[OneHot.scala 58:35]
  assign s2_victim_way = s2_hit_valid ? s2_hit_way : _T_673; // @[DCache.scala 383:26]
  assign releaseWay = _T_2956 ? s2_victim_way : s2_probe_way; // @[DCache.scala 783:81]
  assign _T_321 = inWriteback ? releaseWay : s1_meta_hit_way; // @[DCache.scala 275:61]
  assign _T_332 = {auto_out_d_bits_data[31:24],auto_out_d_bits_data[23:16],auto_out_d_bits_data[15:8],auto_out_d_bits_data[7:0]}; // @[Cat.scala 29:58]
  assign _T_335 = {auto_out_d_bits_data[63:56],auto_out_d_bits_data[55:48],auto_out_d_bits_data[47:40],auto_out_d_bits_data[39:32]}; // @[Cat.scala 29:58]
  assign _T_336 = {auto_out_d_bits_data[63:56],auto_out_d_bits_data[55:48],auto_out_d_bits_data[47:40],auto_out_d_bits_data[39:32],auto_out_d_bits_data[31:24],auto_out_d_bits_data[23:16],auto_out_d_bits_data[15:8],auto_out_d_bits_data[7:0]}; // @[Cat.scala 29:58]
  assign _T_363 = s1_valid_masked & _T_53; // @[DCache.scala 281:28]
  assign _T_367 = &8'hff; // @[DCache.scala 281:93]
  assign _T_368 = ~_T_363 | _T_367; // @[DCache.scala 281:53]
  assign _T_370 = _T_368 | reset; // @[DCache.scala 281:9]
  assign _T_373 = s1_valid_masked & ~s1_sfence; // @[DCache.scala 283:43]
  assign _T_385 = s2_req_cmd == 5'h5; // @[DCache.scala 292:37]
  assign s2_cmd_flush_line = _T_385 & s2_req_size[0]; // @[DCache.scala 293:54]
  assign _T_390 = s1_valid_not_nacked | s1_flush_valid; // @[DCache.scala 297:29]
  assign _T_391_cacheable = tlb_io_resp_cacheable; // @[DCache.scala 301:18]
  assign s2_vaddr = {_T_393[39:12],s2_req_addr[11:0]}; // @[Cat.scala 29:58]
  assign s1_meta_clk_en = _T_390 | s1_probe; // @[DCache.scala 309:62]
  assign s2_meta_corrected_3_tag = _T_465[19:0]; // @[DCache.scala 313:99]
  assign s2_meta_corrected_3_coh_state = _T_465[21:20]; // @[DCache.scala 313:99]
  assign s2_flush_valid = s2_flush_valid_pre_tag_ecc & ~s2_meta_error; // @[DCache.scala 315:51]
  assign _T_471 = s1_valid | inWriteback; // @[DCache.scala 318:23]
  assign en = _T_471 | io_cpu_replay_next; // @[DCache.scala 318:38]
  assign _T_473 = s1_did_read ? 1'h1 : 1'h0; // @[DCache.scala 319:63]
  assign word_en = inWriteback | _T_473; // @[DCache.scala 319:22]
  assign s1_all_data_ways_0 = data_io_resp_0; // @[DCache.scala 277:29 DCache.scala 277:29]
  assign s1_all_data_ways_1 = data_io_resp_1; // @[DCache.scala 277:29 DCache.scala 277:29]
  assign s1_all_data_ways_2 = data_io_resp_2; // @[DCache.scala 277:29 DCache.scala 277:29]
  assign s1_all_data_ways_3 = data_io_resp_3; // @[DCache.scala 277:29 DCache.scala 277:29]
  assign s1_word_en = io_cpu_replay_next ? 1'h1 : word_en; // @[DCache.scala 329:27]
  assign grantIsUncachedData = auto_out_d_bits_opcode == 3'h1; // @[package.scala 15:47]
  assign _T_2877 = blockUncachedGrant | s1_valid; // @[DCache.scala 695:54]
  assign _T_2878 = grantIsUncachedData & _T_2877; // @[DCache.scala 695:31]
  assign grantIsRefill = auto_out_d_bits_opcode == 3'h5; // @[DCache.scala 609:29]
  assign _T_2792 = grantIsRefill & ~dataArb_io_in_1_ready; // @[DCache.scala 665:23]
  assign _T_2745 = auto_out_d_bits_opcode == 3'h4; // @[package.scala 15:47]
  assign grantIsCached = _T_2745 | grantIsRefill; // @[package.scala 64:59]
  assign d_first = _T_2713 == 9'h0; // @[Edges.scala 232:25]
  assign _T_2754 = ~d_first | auto_out_e_ready; // @[DCache.scala 614:50]
  assign canAcceptCachedGrant = ~_T_2956; // @[DCache.scala 613:30]
  assign _T_2755 = _T_2754 & canAcceptCachedGrant; // @[DCache.scala 614:69]
  assign _T_2756 = grantIsCached ? _T_2755 : 1'h1; // @[DCache.scala 614:24]
  assign _GEN_232 = _T_2792 ? 1'h0 : _T_2756; // @[DCache.scala 665:51]
  assign tl_out__d_ready = _T_2878 ? 1'h0 : _GEN_232; // @[DCache.scala 695:68]
  assign _T_2761 = tl_out__d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37]
  assign _T_2722 = auto_out_d_bits_opcode == 3'h0; // @[package.scala 15:47]
  assign _T_2724 = grantIsUncachedData | _T_2722; // @[package.scala 64:59]
  assign _T_2723 = auto_out_d_bits_opcode == 3'h2; // @[package.scala 15:47]
  assign grantIsUncached = _T_2724 | _T_2723; // @[package.scala 64:59]
  assign _GEN_188 = grantIsUncachedData ? 5'h10 : {{1'd0}, _T_321}; // @[DCache.scala 634:34]
  assign _GEN_197 = grantIsUncached ? _GEN_188 : {{1'd0}, _T_321}; // @[DCache.scala 627:35]
  assign _GEN_210 = grantIsCached ? {{1'd0}, _T_321} : _GEN_197; // @[DCache.scala 618:26]
  assign s1_data_way = _T_2761 ? _GEN_210 : {{1'd0}, _T_321}; // @[DCache.scala 617:26]
  assign _T_476 = s1_word_en ? s1_data_way : 5'h0; // @[DCache.scala 331:28]
  assign _T_482 = _T_476[0] ? s1_all_data_ways_0 : 64'h0; // @[Mux.scala 27:72]
  assign _T_483 = _T_476[1] ? s1_all_data_ways_1 : 64'h0; // @[Mux.scala 27:72]
  assign _T_484 = _T_476[2] ? s1_all_data_ways_2 : 64'h0; // @[Mux.scala 27:72]
  assign _T_485 = _T_476[3] ? s1_all_data_ways_3 : 64'h0; // @[Mux.scala 27:72]
  assign _T_486 = _T_476[4] ? _T_336 : 64'h0; // @[Mux.scala 27:72]
  assign _T_487 = _T_482 | _T_483; // @[Mux.scala 27:72]
  assign _T_488 = _T_487 | _T_484; // @[Mux.scala 27:72]
  assign _T_489 = _T_488 | _T_485; // @[Mux.scala 27:72]
  assign _T_490 = _T_489 | _T_486; // @[Mux.scala 27:72]
  assign _T_633 = {s2_data[31:24],s2_data[23:16],s2_data[15:8],s2_data[7:0]}; // @[Cat.scala 29:58]
  assign _T_636 = {s2_data[63:56],s2_data[55:48],s2_data[47:40],s2_data[39:32]}; // @[Cat.scala 29:58]
  assign s2_data_corrected = {s2_data[63:56],s2_data[55:48],s2_data[47:40],s2_data[39:32],s2_data[31:24],s2_data[23:16],s2_data[15:8],s2_data[7:0]}; // @[Cat.scala 29:58]
  assign s2_valid_flush_line = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_cmd_flush_line; // @[DCache.scala 371:75]
  assign _T_650 = s2_valid_masked & s2_readwrite; // @[DCache.scala 375:39]
  assign _T_652 = _T_650 & ~s2_meta_error; // @[DCache.scala 375:55]
  assign s2_valid_miss = _T_652 & ~s2_hit; // @[DCache.scala 375:73]
  assign s2_uncached = ~s2_pma_cacheable; // @[DCache.scala 376:21]
  assign _T_660 = s2_valid_miss & ~s2_uncached; // @[DCache.scala 377:44]
  assign _T_661 = |uncachedInFlight_0; // @[DCache.scala 377:88]
  assign s2_valid_cached_miss = _T_660 & ~_T_661; // @[DCache.scala 377:60]
  assign _T_663 = s2_valid_cached_miss | s2_valid_flush_line; // @[DCache.scala 379:79]
  assign s2_want_victimize = _T_663 | s2_flush_valid; // @[DCache.scala 379:125]
  assign _T_668 = s2_valid_miss & s2_uncached; // @[DCache.scala 382:49]
  assign _T_669 = &uncachedInFlight_0; // @[DCache.scala 382:92]
  assign s2_valid_uncached_pending = _T_668 & ~_T_669; // @[DCache.scala 382:64]
  assign s2_victim_tag = s2_valid_flush_line ? s2_req_addr[31:12] : _T_677; // @[DCache.scala 384:26]
  assign s2_victim_state_state = s2_hit_valid ? s2_hit_state_state : _T_679_state; // @[DCache.scala 385:28]
  assign _T_695 = _T_693 ? 3'h5 : 3'h0; // @[Misc.scala 37:36]
  assign _T_699 = _T_697 ? 3'h2 : _T_695; // @[Misc.scala 37:36]
  assign _T_703 = _T_701 ? 3'h1 : _T_699; // @[Misc.scala 37:36]
  assign _T_707 = _T_705 ? 3'h1 : _T_703; // @[Misc.scala 37:36]
  assign _T_711 = _T_709 ? 3'h5 : _T_707; // @[Misc.scala 37:36]
  assign _T_715 = _T_713 ? 3'h4 : _T_711; // @[Misc.scala 37:36]
  assign _T_716 = _T_713 ? 2'h1 : 2'h0; // @[Misc.scala 37:63]
  assign _T_719 = _T_717 ? 3'h0 : _T_715; // @[Misc.scala 37:36]
  assign _T_720 = _T_717 ? 2'h1 : _T_716; // @[Misc.scala 37:63]
  assign _T_723 = _T_721 ? 3'h0 : _T_719; // @[Misc.scala 37:36]
  assign _T_724 = _T_721 ? 2'h1 : _T_720; // @[Misc.scala 37:63]
  assign _T_727 = _T_725 ? 3'h5 : _T_723; // @[Misc.scala 37:36]
  assign _T_728 = _T_725 ? 2'h0 : _T_724; // @[Misc.scala 37:63]
  assign _T_731 = _T_729 ? 3'h4 : _T_727; // @[Misc.scala 37:36]
  assign _T_732 = _T_729 ? 2'h1 : _T_728; // @[Misc.scala 37:63]
  assign _T_735 = _T_733 ? 3'h3 : _T_731; // @[Misc.scala 37:36]
  assign _T_736 = _T_733 ? 2'h2 : _T_732; // @[Misc.scala 37:63]
  assign s2_report_param = _T_737 ? 3'h3 : _T_735; // @[Misc.scala 37:36]
  assign probeNewCoh_state = _T_737 ? 2'h2 : _T_736; // @[Misc.scala 37:63]
  assign _T_745 = {2'h2,s2_victim_state_state}; // @[Cat.scala 29:58]
  assign _T_758 = 4'h8 == _T_745; // @[Misc.scala 55:20]
  assign _T_760 = _T_758 ? 3'h5 : 3'h0; // @[Misc.scala 37:36]
  assign _T_762 = 4'h9 == _T_745; // @[Misc.scala 55:20]
  assign _T_764 = _T_762 ? 3'h2 : _T_760; // @[Misc.scala 37:36]
  assign _T_766 = 4'ha == _T_745; // @[Misc.scala 55:20]
  assign _T_768 = _T_766 ? 3'h1 : _T_764; // @[Misc.scala 37:36]
  assign _T_770 = 4'hb == _T_745; // @[Misc.scala 55:20]
  assign _T_772 = _T_770 ? 3'h1 : _T_768; // @[Misc.scala 37:36]
  assign _T_774 = 4'h4 == _T_745; // @[Misc.scala 55:20]
  assign _T_775 = _T_774 ? 1'h0 : _T_770; // @[Misc.scala 37:9]
  assign _T_776 = _T_774 ? 3'h5 : _T_772; // @[Misc.scala 37:36]
  assign _T_778 = 4'h5 == _T_745; // @[Misc.scala 55:20]
  assign _T_779 = _T_778 ? 1'h0 : _T_775; // @[Misc.scala 37:9]
  assign _T_780 = _T_778 ? 3'h4 : _T_776; // @[Misc.scala 37:36]
  assign _T_781 = _T_778 ? 2'h1 : 2'h0; // @[Misc.scala 37:63]
  assign _T_782 = 4'h6 == _T_745; // @[Misc.scala 55:20]
  assign _T_783 = _T_782 ? 1'h0 : _T_779; // @[Misc.scala 37:9]
  assign _T_784 = _T_782 ? 3'h0 : _T_780; // @[Misc.scala 37:36]
  assign _T_785 = _T_782 ? 2'h1 : _T_781; // @[Misc.scala 37:63]
  assign _T_786 = 4'h7 == _T_745; // @[Misc.scala 55:20]
  assign _T_787 = _T_786 | _T_783; // @[Misc.scala 37:9]
  assign _T_788 = _T_786 ? 3'h0 : _T_784; // @[Misc.scala 37:36]
  assign _T_789 = _T_786 ? 2'h1 : _T_785; // @[Misc.scala 37:63]
  assign _T_790 = 4'h0 == _T_745; // @[Misc.scala 55:20]
  assign _T_791 = _T_790 ? 1'h0 : _T_787; // @[Misc.scala 37:9]
  assign _T_792 = _T_790 ? 3'h5 : _T_788; // @[Misc.scala 37:36]
  assign _T_793 = _T_790 ? 2'h0 : _T_789; // @[Misc.scala 37:63]
  assign _T_794 = 4'h1 == _T_745; // @[Misc.scala 55:20]
  assign _T_795 = _T_794 ? 1'h0 : _T_791; // @[Misc.scala 37:9]
  assign _T_796 = _T_794 ? 3'h4 : _T_792; // @[Misc.scala 37:36]
  assign _T_797 = _T_794 ? 2'h1 : _T_793; // @[Misc.scala 37:63]
  assign _T_798 = 4'h2 == _T_745; // @[Misc.scala 55:20]
  assign _T_799 = _T_798 ? 1'h0 : _T_795; // @[Misc.scala 37:9]
  assign _T_800 = _T_798 ? 3'h3 : _T_796; // @[Misc.scala 37:36]
  assign _T_801 = _T_798 ? 2'h2 : _T_797; // @[Misc.scala 37:63]
  assign _T_802 = 4'h3 == _T_745; // @[Misc.scala 55:20]
  assign s2_victim_dirty = _T_802 | _T_799; // @[Misc.scala 37:9]
  assign s2_shrink_param = _T_802 ? 3'h3 : _T_800; // @[Misc.scala 37:36]
  assign voluntaryNewCoh_state = _T_802 ? 2'h2 : _T_801; // @[Misc.scala 37:63]
  assign s2_dont_nack_uncached = s2_valid_uncached_pending & auto_out_a_ready; // @[DCache.scala 391:57]
  assign _T_815 = s2_req_cmd == 5'h17; // @[DCache.scala 395:17]
  assign s2_dont_nack_misc = _T_644 & _T_815; // @[DCache.scala 392:61]
  assign _T_818 = s2_valid_no_xcpt & ~s2_dont_nack_uncached; // @[DCache.scala 396:38]
  assign _T_820 = _T_818 & ~s2_dont_nack_misc; // @[DCache.scala 396:64]
  assign _T_831 = s2_valid_masked | s2_flush_valid_pre_tag_ecc; // @[DCache.scala 401:63]
  assign _T_832 = _T_831 | s2_probe; // @[DCache.scala 401:93]
  assign _T_848 = {metaArb_io_in_1_bits_idx, 6'h0}; // @[DCache.scala 405:98]
  assign new_meta_coh_state = s2_meta_error ? 2'h0 : s2_meta_corrected_3_coh_state; // @[DCache.scala 408:40]
  assign _T_863 = lrscCount > 7'h0; // @[DCache.scala 425:34]
  assign lrscBackingOff = _T_863 & ~lrscValid; // @[DCache.scala 425:38]
  assign lrscAddrMatch = lrscAddr == s2_req_addr[39:6]; // @[DCache.scala 427:32]
  assign _T_866 = lrscValid & lrscAddrMatch; // @[DCache.scala 428:41]
  assign s2_sc_fail = _T_421 & ~_T_866; // @[DCache.scala 428:26]
  assign _T_868 = s2_valid_hit_pre_data_ecc_and_waw & _T_541; // @[DCache.scala 429:23]
  assign _T_870 = _T_868 & ~cached_grant_wait; // @[DCache.scala 429:32]
  assign _T_871 = _T_870 | s2_valid_cached_miss; // @[DCache.scala 429:54]
  assign _T_878 = lrscCount - 7'h1; // @[DCache.scala 433:49]
  assign _T_879 = s2_valid_masked & lrscValid; // @[DCache.scala 434:29]
  assign _T_887 = s1_valid_not_nacked & s1_write; // @[DCache.scala 443:63]
  assign _T_941 = s1_write & _T_53; // @[DCache.scala 1086:23]
  assign _T_942 = s1_read | _T_941; // @[DCache.scala 1085:21]
  assign _T_946 = s2_valid_hit_pre_data_ecc_and_waw & s2_write; // @[DCache.scala 441:46]
  assign _T_948 = _T_946 & ~s2_sc_fail; // @[DCache.scala 441:58]
  assign pstore_drain_opportunistic = ~_T_167; // @[DCache.scala 453:36]
  assign pstore_drain_on_miss = releaseInFlight | _T_1016; // @[DCache.scala 454:46]
  assign pstore1_valid = _T_948 | pstore1_held; // @[DCache.scala 458:38]
  assign _T_1024 = pstore1_valid_likely & pstore2_valid; // @[DCache.scala 460:54]
  assign _T_1025 = s1_valid & s1_write; // @[DCache.scala 460:85]
  assign _T_1026 = _T_1025 | pstore1_rmw; // @[DCache.scala 460:98]
  assign pstore_drain_structural = _T_1024 & _T_1026; // @[DCache.scala 460:71]
  assign _T_1030 = _T_946 | pstore1_held; // @[DCache.scala 457:96]
  assign _T_1031 = _T_1030 == pstore1_valid; // @[DCache.scala 461:63]
  assign _T_1032 = pstore1_rmw | _T_1031; // @[DCache.scala 461:22]
  assign _T_1034 = _T_1032 | reset; // @[DCache.scala 461:9]
  assign _T_1045 = _T_1030 & ~pstore1_rmw; // @[DCache.scala 469:41]
  assign _T_1046 = _T_1045 | pstore2_valid; // @[DCache.scala 469:58]
  assign _T_1047 = pstore_drain_opportunistic | pstore_drain_on_miss; // @[DCache.scala 469:107]
  assign _T_1048 = _T_1046 & _T_1047; // @[DCache.scala 469:76]
  assign pstore_drain = pstore_drain_structural | _T_1048; // @[DCache.scala 468:48]
  assign _T_1058 = pstore1_valid & pstore2_valid; // @[DCache.scala 472:71]
  assign _T_1062 = pstore2_valid == pstore_drain; // @[DCache.scala 473:79]
  assign advance_pstore1 = pstore1_valid & _T_1062; // @[DCache.scala 473:61]
  assign _T_1064 = pstore2_valid & ~pstore_drain; // @[DCache.scala 474:34]
  assign pstore1_storegen_data = amoalu_io_out; // @[DCache.scala 888:27]
  assign pstore2_storegen_data = {_T_1107,_T_1102,_T_1097,_T_1092,_T_1087,_T_1082,_T_1077,_T_1072}; // @[Cat.scala 29:58]
  assign _T_1132 = pstore2_valid ? pstore2_addr : pstore1_addr; // @[DCache.scala 500:36]
  assign _T_1134 = pstore2_valid ? pstore2_storegen_data : pstore1_data; // @[DCache.scala 502:63]
  assign _T_1145 = {_T_1134[31:24],_T_1134[23:16],_T_1134[15:8],_T_1134[7:0]}; // @[Cat.scala 29:58]
  assign _T_1148 = {_T_1134[63:56],_T_1134[55:48],_T_1134[47:40],_T_1134[39:32]}; // @[Cat.scala 29:58]
  assign _T_1152 = pstore2_valid ? mask : pstore1_mask; // @[DCache.scala 504:47]
  assign _T_1161 = |_T_1152[0]; // @[DCache.scala 1076:66]
  assign _T_1162 = |_T_1152[1]; // @[DCache.scala 1076:66]
  assign _T_1163 = |_T_1152[2]; // @[DCache.scala 1076:66]
  assign _T_1164 = |_T_1152[3]; // @[DCache.scala 1076:66]
  assign _T_1165 = |_T_1152[4]; // @[DCache.scala 1076:66]
  assign _T_1166 = |_T_1152[5]; // @[DCache.scala 1076:66]
  assign _T_1167 = |_T_1152[6]; // @[DCache.scala 1076:66]
  assign _T_1168 = |_T_1152[7]; // @[DCache.scala 1076:66]
  assign _T_1171 = {_T_1164,_T_1163,_T_1162,_T_1161}; // @[Cat.scala 29:58]
  assign _T_1174 = {_T_1168,_T_1167,_T_1166,_T_1165}; // @[Cat.scala 29:58]
  assign _T_1355 = {~uncachedInFlight_0, 1'h0}; // @[DCache.scala 524:59]
  assign a_source = _T_1355[0] ? 1'h0 : 1'h1; // @[Mux.scala 47:69]
  assign acquire_address = {s2_req_addr[39:6], 6'h0}; // @[DCache.scala 525:49]
  assign a_mask = {{15'd0}, pstore1_mask}; // @[DCache.scala 529:29]
  assign _T_1412 = {{1'd0}, s2_req_size}; // @[Misc.scala 201:34]
  assign _T_1414 = 4'h1 << _T_1412[1:0]; // @[OneHot.scala 65:12]
  assign _T_1416 = _T_1414[2:0] | 3'h1; // @[Misc.scala 201:81]
  assign _T_1417 = s2_req_size >= 2'h3; // @[Misc.scala 205:21]
  assign _T_1422 = _T_1416[2] & ~s2_req_addr[2]; // @[Misc.scala 214:38]
  assign _T_1423 = _T_1417 | _T_1422; // @[Misc.scala 214:29]
  assign _T_1425 = _T_1416[2] & s2_req_addr[2]; // @[Misc.scala 214:38]
  assign _T_1426 = _T_1417 | _T_1425; // @[Misc.scala 214:29]
  assign _T_1430 = ~s2_req_addr[2] & ~s2_req_addr[1]; // @[Misc.scala 213:27]
  assign _T_1431 = _T_1416[1] & _T_1430; // @[Misc.scala 214:38]
  assign _T_1432 = _T_1423 | _T_1431; // @[Misc.scala 214:29]
  assign _T_1433 = ~s2_req_addr[2] & s2_req_addr[1]; // @[Misc.scala 213:27]
  assign _T_1434 = _T_1416[1] & _T_1433; // @[Misc.scala 214:38]
  assign _T_1435 = _T_1423 | _T_1434; // @[Misc.scala 214:29]
  assign _T_1436 = s2_req_addr[2] & ~s2_req_addr[1]; // @[Misc.scala 213:27]
  assign _T_1437 = _T_1416[1] & _T_1436; // @[Misc.scala 214:38]
  assign _T_1438 = _T_1426 | _T_1437; // @[Misc.scala 214:29]
  assign _T_1439 = s2_req_addr[2] & s2_req_addr[1]; // @[Misc.scala 213:27]
  assign _T_1440 = _T_1416[1] & _T_1439; // @[Misc.scala 214:38]
  assign _T_1441 = _T_1426 | _T_1440; // @[Misc.scala 214:29]
  assign _T_1445 = _T_1430 & ~s2_req_addr[0]; // @[Misc.scala 213:27]
  assign _T_1446 = _T_1416[0] & _T_1445; // @[Misc.scala 214:38]
  assign _T_1447 = _T_1432 | _T_1446; // @[Misc.scala 214:29]
  assign _T_1448 = _T_1430 & s2_req_addr[0]; // @[Misc.scala 213:27]
  assign _T_1449 = _T_1416[0] & _T_1448; // @[Misc.scala 214:38]
  assign _T_1450 = _T_1432 | _T_1449; // @[Misc.scala 214:29]
  assign _T_1451 = _T_1433 & ~s2_req_addr[0]; // @[Misc.scala 213:27]
  assign _T_1452 = _T_1416[0] & _T_1451; // @[Misc.scala 214:38]
  assign _T_1453 = _T_1435 | _T_1452; // @[Misc.scala 214:29]
  assign _T_1454 = _T_1433 & s2_req_addr[0]; // @[Misc.scala 213:27]
  assign _T_1455 = _T_1416[0] & _T_1454; // @[Misc.scala 214:38]
  assign _T_1456 = _T_1435 | _T_1455; // @[Misc.scala 214:29]
  assign _T_1457 = _T_1436 & ~s2_req_addr[0]; // @[Misc.scala 213:27]
  assign _T_1458 = _T_1416[0] & _T_1457; // @[Misc.scala 214:38]
  assign _T_1459 = _T_1438 | _T_1458; // @[Misc.scala 214:29]
  assign _T_1460 = _T_1436 & s2_req_addr[0]; // @[Misc.scala 213:27]
  assign _T_1461 = _T_1416[0] & _T_1460; // @[Misc.scala 214:38]
  assign _T_1462 = _T_1438 | _T_1461; // @[Misc.scala 214:29]
  assign _T_1463 = _T_1439 & ~s2_req_addr[0]; // @[Misc.scala 213:27]
  assign _T_1464 = _T_1416[0] & _T_1463; // @[Misc.scala 214:38]
  assign _T_1465 = _T_1441 | _T_1464; // @[Misc.scala 214:29]
  assign _T_1466 = _T_1439 & s2_req_addr[0]; // @[Misc.scala 213:27]
  assign _T_1467 = _T_1416[0] & _T_1466; // @[Misc.scala 214:38]
  assign _T_1468 = _T_1441 | _T_1467; // @[Misc.scala 214:29]
  assign get_mask = {_T_1468,_T_1465,_T_1462,_T_1459,_T_1456,_T_1453,_T_1450,_T_1447}; // @[Cat.scala 29:58]
  assign _T_2577 = 5'h4 == s2_req_cmd; // @[Mux.scala 80:60]
  assign _T_2578_opcode = _T_2577 ? 3'h3 : 3'h0; // @[Mux.scala 80:57]
  assign _T_1696_size = {{2'd0}, s2_req_size}; // @[Edges.scala 515:17 Edges.scala 518:15]
  assign _T_2578_size = _T_2577 ? _T_1696_size : 4'h0; // @[Mux.scala 80:57]
  assign _T_2578_source = _T_2577 & a_source; // @[Mux.scala 80:57]
  assign _T_2578_address = _T_2577 ? s2_req_addr[31:0] : 32'h0; // @[Mux.scala 80:57]
  assign _T_2578_mask = _T_2577 ? get_mask : 8'h0; // @[Mux.scala 80:57]
  assign _T_2578_data = _T_2577 ? pstore1_data : 64'h0; // @[Mux.scala 80:57]
  assign _T_2579 = 5'h9 == s2_req_cmd; // @[Mux.scala 80:60]
  assign _T_2580_opcode = _T_2579 ? 3'h3 : _T_2578_opcode; // @[Mux.scala 80:57]
  assign _T_2580_param = _T_2579 ? 3'h0 : _T_2578_opcode; // @[Mux.scala 80:57]
  assign _T_2580_size = _T_2579 ? _T_1696_size : _T_2578_size; // @[Mux.scala 80:57]
  assign _T_2580_source = _T_2579 ? a_source : _T_2578_source; // @[Mux.scala 80:57]
  assign _T_2580_address = _T_2579 ? s2_req_addr[31:0] : _T_2578_address; // @[Mux.scala 80:57]
  assign _T_2580_mask = _T_2579 ? get_mask : _T_2578_mask; // @[Mux.scala 80:57]
  assign _T_2580_data = _T_2579 ? pstore1_data : _T_2578_data; // @[Mux.scala 80:57]
  assign _T_2581 = 5'ha == s2_req_cmd; // @[Mux.scala 80:60]
  assign _T_2582_opcode = _T_2581 ? 3'h3 : _T_2580_opcode; // @[Mux.scala 80:57]
  assign _T_2582_param = _T_2581 ? 3'h1 : _T_2580_param; // @[Mux.scala 80:57]
  assign _T_2582_size = _T_2581 ? _T_1696_size : _T_2580_size; // @[Mux.scala 80:57]
  assign _T_2582_source = _T_2581 ? a_source : _T_2580_source; // @[Mux.scala 80:57]
  assign _T_2582_address = _T_2581 ? s2_req_addr[31:0] : _T_2580_address; // @[Mux.scala 80:57]
  assign _T_2582_mask = _T_2581 ? get_mask : _T_2580_mask; // @[Mux.scala 80:57]
  assign _T_2582_data = _T_2581 ? pstore1_data : _T_2580_data; // @[Mux.scala 80:57]
  assign _T_2583 = 5'hb == s2_req_cmd; // @[Mux.scala 80:60]
  assign _T_2584_opcode = _T_2583 ? 3'h3 : _T_2582_opcode; // @[Mux.scala 80:57]
  assign _T_2584_param = _T_2583 ? 3'h2 : _T_2582_param; // @[Mux.scala 80:57]
  assign _T_2584_size = _T_2583 ? _T_1696_size : _T_2582_size; // @[Mux.scala 80:57]
  assign _T_2584_source = _T_2583 ? a_source : _T_2582_source; // @[Mux.scala 80:57]
  assign _T_2584_address = _T_2583 ? s2_req_addr[31:0] : _T_2582_address; // @[Mux.scala 80:57]
  assign _T_2584_mask = _T_2583 ? get_mask : _T_2582_mask; // @[Mux.scala 80:57]
  assign _T_2584_data = _T_2583 ? pstore1_data : _T_2582_data; // @[Mux.scala 80:57]
  assign _T_2585 = 5'h8 == s2_req_cmd; // @[Mux.scala 80:60]
  assign _T_2586_opcode = _T_2585 ? 3'h2 : _T_2584_opcode; // @[Mux.scala 80:57]
  assign _T_2586_param = _T_2585 ? 3'h4 : _T_2584_param; // @[Mux.scala 80:57]
  assign _T_2586_size = _T_2585 ? _T_1696_size : _T_2584_size; // @[Mux.scala 80:57]
  assign _T_2586_source = _T_2585 ? a_source : _T_2584_source; // @[Mux.scala 80:57]
  assign _T_2586_address = _T_2585 ? s2_req_addr[31:0] : _T_2584_address; // @[Mux.scala 80:57]
  assign _T_2586_mask = _T_2585 ? get_mask : _T_2584_mask; // @[Mux.scala 80:57]
  assign _T_2586_data = _T_2585 ? pstore1_data : _T_2584_data; // @[Mux.scala 80:57]
  assign _T_2587 = 5'hc == s2_req_cmd; // @[Mux.scala 80:60]
  assign _T_2588_opcode = _T_2587 ? 3'h2 : _T_2586_opcode; // @[Mux.scala 80:57]
  assign _T_2588_param = _T_2587 ? 3'h0 : _T_2586_param; // @[Mux.scala 80:57]
  assign _T_2588_size = _T_2587 ? _T_1696_size : _T_2586_size; // @[Mux.scala 80:57]
  assign _T_2588_source = _T_2587 ? a_source : _T_2586_source; // @[Mux.scala 80:57]
  assign _T_2588_address = _T_2587 ? s2_req_addr[31:0] : _T_2586_address; // @[Mux.scala 80:57]
  assign _T_2588_mask = _T_2587 ? get_mask : _T_2586_mask; // @[Mux.scala 80:57]
  assign _T_2588_data = _T_2587 ? pstore1_data : _T_2586_data; // @[Mux.scala 80:57]
  assign _T_2589 = 5'hd == s2_req_cmd; // @[Mux.scala 80:60]
  assign _T_2590_opcode = _T_2589 ? 3'h2 : _T_2588_opcode; // @[Mux.scala 80:57]
  assign _T_2590_param = _T_2589 ? 3'h1 : _T_2588_param; // @[Mux.scala 80:57]
  assign _T_2590_size = _T_2589 ? _T_1696_size : _T_2588_size; // @[Mux.scala 80:57]
  assign _T_2590_source = _T_2589 ? a_source : _T_2588_source; // @[Mux.scala 80:57]
  assign _T_2590_address = _T_2589 ? s2_req_addr[31:0] : _T_2588_address; // @[Mux.scala 80:57]
  assign _T_2590_mask = _T_2589 ? get_mask : _T_2588_mask; // @[Mux.scala 80:57]
  assign _T_2590_data = _T_2589 ? pstore1_data : _T_2588_data; // @[Mux.scala 80:57]
  assign _T_2591 = 5'he == s2_req_cmd; // @[Mux.scala 80:60]
  assign _T_2592_opcode = _T_2591 ? 3'h2 : _T_2590_opcode; // @[Mux.scala 80:57]
  assign _T_2592_param = _T_2591 ? 3'h2 : _T_2590_param; // @[Mux.scala 80:57]
  assign _T_2592_size = _T_2591 ? _T_1696_size : _T_2590_size; // @[Mux.scala 80:57]
  assign _T_2592_source = _T_2591 ? a_source : _T_2590_source; // @[Mux.scala 80:57]
  assign _T_2592_address = _T_2591 ? s2_req_addr[31:0] : _T_2590_address; // @[Mux.scala 80:57]
  assign _T_2592_mask = _T_2591 ? get_mask : _T_2590_mask; // @[Mux.scala 80:57]
  assign _T_2592_data = _T_2591 ? pstore1_data : _T_2590_data; // @[Mux.scala 80:57]
  assign _T_2593 = 5'hf == s2_req_cmd; // @[Mux.scala 80:60]
  assign atomics_opcode = _T_2593 ? 3'h2 : _T_2592_opcode; // @[Mux.scala 80:57]
  assign atomics_param = _T_2593 ? 3'h3 : _T_2592_param; // @[Mux.scala 80:57]
  assign atomics_size = _T_2593 ? _T_1696_size : _T_2592_size; // @[Mux.scala 80:57]
  assign atomics_source = _T_2593 ? a_source : _T_2592_source; // @[Mux.scala 80:57]
  assign atomics_address = _T_2593 ? s2_req_addr[31:0] : _T_2592_address; // @[Mux.scala 80:57]
  assign atomics_mask = _T_2593 ? get_mask : _T_2592_mask; // @[Mux.scala 80:57]
  assign atomics_data = _T_2593 ? pstore1_data : _T_2592_data; // @[Mux.scala 80:57]
  assign _T_2596 = s2_valid_cached_miss & ~release_ack_wait; // @[DCache.scala 551:27]
  assign _T_2600 = _T_2596 & ~s2_victim_dirty; // @[DCache.scala 551:48]
  assign tl_out_a_valid = s2_valid_uncached_pending | _T_2600; // @[DCache.scala 550:67]
  assign _T_2693_opcode = s2_read ? atomics_opcode : 3'h0; // @[DCache.scala 555:8]
  assign _T_2693_param = s2_read ? atomics_param : 3'h0; // @[DCache.scala 555:8]
  assign _T_2693_size = s2_read ? atomics_size : _T_1696_size; // @[DCache.scala 555:8]
  assign _T_2693_source = s2_read ? atomics_source : a_source; // @[DCache.scala 555:8]
  assign _T_2693_address = s2_read ? atomics_address : s2_req_addr[31:0]; // @[DCache.scala 555:8]
  assign _T_2693_mask = s2_read ? atomics_mask : get_mask; // @[DCache.scala 555:8]
  assign _T_2693_data = s2_read ? atomics_data : pstore1_data; // @[DCache.scala 555:8]
  assign _T_2694_opcode = _T_419 ? 3'h1 : _T_2693_opcode; // @[DCache.scala 554:8]
  assign _T_2694_param = _T_419 ? 3'h0 : _T_2693_param; // @[DCache.scala 554:8]
  assign _T_2694_size = _T_419 ? _T_1696_size : _T_2693_size; // @[DCache.scala 554:8]
  assign _T_2694_source = _T_419 ? a_source : _T_2693_source; // @[DCache.scala 554:8]
  assign _T_2694_address = _T_419 ? s2_req_addr[31:0] : _T_2693_address; // @[DCache.scala 554:8]
  assign putpartial_mask = a_mask[7:0]; // @[Edges.scala 485:17 Edges.scala 491:15]
  assign _T_2694_mask = _T_419 ? putpartial_mask : _T_2693_mask; // @[DCache.scala 554:8]
  assign _T_2694_data = _T_419 ? pstore1_data : _T_2693_data; // @[DCache.scala 554:8]
  assign _T_2695_opcode = s2_write ? _T_2694_opcode : 3'h4; // @[DCache.scala 553:8]
  assign _T_2695_param = s2_write ? _T_2694_param : 3'h0; // @[DCache.scala 553:8]
  assign _T_2695_size = s2_write ? _T_2694_size : _T_1696_size; // @[DCache.scala 553:8]
  assign _T_2695_source = s2_write ? _T_2694_source : a_source; // @[DCache.scala 553:8]
  assign _T_2695_address = s2_write ? _T_2694_address : s2_req_addr[31:0]; // @[DCache.scala 553:8]
  assign _T_2695_mask = s2_write ? _T_2694_mask : get_mask; // @[DCache.scala 553:8]
  assign _T_2695_data = s2_write ? _T_2694_data : 64'h0; // @[DCache.scala 553:8]
  assign _T_2625_param = {{1'd0}, s2_grow_param}; // @[Edges.scala 347:17 Edges.scala 349:15]
  assign _T_2698 = 2'h1 << a_source; // @[OneHot.scala 65:12]
  assign a_sel = _T_2698[1]; // @[DCache.scala 574:66]
  assign _T_2700 = auto_out_a_ready & tl_out_a_valid; // @[Decoupled.scala 40:37]
  assign _GEN_143 = a_sel | uncachedInFlight_0; // @[DCache.scala 578:18]
  assign _T_2707 = 27'hfff << auto_out_d_bits_size; // @[package.scala 212:77]
  assign _T_2710 = ~_T_2707[11:3]; // @[Edges.scala 221:59]
  assign _T_2712 = auto_out_d_bits_opcode[0] ? _T_2710 : 9'h0; // @[Edges.scala 222:14]
  assign _T_2715 = _T_2713 - 9'h1; // @[Edges.scala 231:28]
  assign _T_2716 = _T_2713 == 9'h1; // @[Edges.scala 233:25]
  assign _T_2717 = _T_2712 == 9'h0; // @[Edges.scala 233:47]
  assign d_last = _T_2716 | _T_2717; // @[Edges.scala 233:37]
  assign d_done = d_last & _T_2761; // @[Edges.scala 234:22]
  assign _T_2719 = _T_2712 & ~_T_2715; // @[Edges.scala 235:25]
  assign d_address_inc = {_T_2719, 3'h0}; // @[Edges.scala 270:29]
  assign grantIsVoluntary = auto_out_d_bits_opcode == 3'h6; // @[DCache.scala 608:32]
  assign _T_2749 = blockProbeAfterGrantCount - 3'h1; // @[DCache.scala 612:97]
  assign _T_2758 = 2'h1 << auto_out_d_bits_source; // @[OneHot.scala 65:12]
  assign uncachedRespIdxOH = _T_2758[1]; // @[DCache.scala 615:90]
  assign _T_2763 = cached_grant_wait | reset; // @[DCache.scala 620:13]
  assign _T_2766 = uncachedRespIdxOH & d_last; // @[DCache.scala 629:17]
  assign _T_2768 = uncachedInFlight_0 | reset; // @[DCache.scala 630:17]
  assign dontCareBits = {s1_paddr[31:3], 3'h0}; // @[DCache.scala 644:55]
  assign _GEN_347 = {{29'd0}, uncachedReqs_0_addr[2:0]}; // @[DCache.scala 645:26]
  assign _T_2773 = dontCareBits | _GEN_347; // @[DCache.scala 645:26]
  assign _T_2775 = release_ack_wait | reset; // @[DCache.scala 651:13]
  assign _GEN_195 = grantIsVoluntary ? 1'h0 : release_ack_wait; // @[DCache.scala 650:36]
  assign _GEN_204 = grantIsUncached ? release_ack_wait : _GEN_195; // @[DCache.scala 627:35]
  assign _GEN_208 = grantIsCached & d_last; // @[DCache.scala 618:26]
  assign _GEN_217 = grantIsCached ? release_ack_wait : _GEN_204; // @[DCache.scala 618:26]
  assign _GEN_230 = _T_2761 ? _GEN_217 : release_ack_wait; // @[DCache.scala 617:26]
  assign _T_2777 = auto_out_d_valid & d_first; // @[DCache.scala 657:36]
  assign _T_2778 = _T_2777 & grantIsCached; // @[DCache.scala 657:47]
  assign _T_2779 = _T_2778 & canAcceptCachedGrant; // @[DCache.scala 657:64]
  assign tl_out__e_valid = _T_2792 ? 1'h0 : _T_2779; // @[DCache.scala 665:51]
  assign _T_2781 = auto_out_e_ready & tl_out__e_valid; // @[Decoupled.scala 40:37]
  assign _T_2783 = _T_2761 & d_first; // @[DCache.scala 659:47]
  assign _T_2784 = _T_2783 & grantIsCached; // @[DCache.scala 659:58]
  assign _T_2785 = _T_2781 == _T_2784; // @[DCache.scala 659:26]
  assign _T_2787 = _T_2785 | reset; // @[DCache.scala 659:9]
  assign _T_2789 = auto_out_d_valid & grantIsRefill; // @[DCache.scala 664:44]
  assign _T_2790 = _T_2789 & canAcceptCachedGrant; // @[DCache.scala 664:61]
  assign _T_2794 = {s2_vaddr[39:6], 6'h0}; // @[DCache.scala 671:57]
  assign _GEN_348 = {{28'd0}, d_address_inc}; // @[DCache.scala 671:67]
  assign _T_2795 = _T_2794 | _GEN_348; // @[DCache.scala 671:67]
  assign _T_2798 = grantIsCached & d_done; // @[DCache.scala 684:43]
  assign _T_2857 = {s2_write,_T_542,auto_out_d_bits_param}; // @[Cat.scala 29:58]
  assign _T_2866 = 4'h1 == _T_2857; // @[Mux.scala 80:60]
  assign _T_2867 = _T_2866 ? 2'h1 : 2'h0; // @[Mux.scala 80:57]
  assign _T_2868 = 4'h0 == _T_2857; // @[Mux.scala 80:60]
  assign _T_2869 = _T_2868 ? 2'h2 : _T_2867; // @[Mux.scala 80:57]
  assign _T_2870 = 4'h4 == _T_2857; // @[Mux.scala 80:60]
  assign _T_2871 = _T_2870 ? 2'h2 : _T_2869; // @[Mux.scala 80:57]
  assign _T_2872 = 4'hc == _T_2857; // @[Mux.scala 80:60]
  assign _T_2873 = _T_2872 ? 2'h3 : _T_2871; // @[Mux.scala 80:57]
  assign _GEN_233 = auto_out_d_valid ? 1'h0 : _GEN_31; // @[DCache.scala 698:29]
  assign _GEN_234 = auto_out_d_valid | _T_2790; // @[DCache.scala 698:29]
  assign _GEN_235 = auto_out_d_valid ? 1'h0 : 1'h1; // @[DCache.scala 698:29]
  assign _T_2888 = ~block_probe_for_core_progress | lrscBackingOff; // @[DCache.scala 712:79]
  assign _T_2889 = auto_out_b_valid & _T_2888; // @[DCache.scala 712:44]
  assign _T_2897 = {io_cpu_req_bits_addr[39:32],auto_out_b_bits_address}; // @[Cat.scala 29:58]
  assign _T_2908 = _T_2906 - 9'h1; // @[Edges.scala 231:28]
  assign c_count = _T_2905 & ~_T_2908; // @[Edges.scala 235:25]
  assign releaseRejected = s2_release_data_valid & ~_T_2898; // @[DCache.scala 725:44]
  assign _T_2919 = {1'h0,c_count}; // @[Cat.scala 29:58]
  assign _T_2920 = {1'h0,s2_release_data_valid}; // @[Cat.scala 29:58]
  assign _GEN_349 = {{1'd0}, s1_release_data_valid}; // @[DCache.scala 726:101]
  assign _T_2922 = _GEN_349 + _T_2920; // @[DCache.scala 726:101]
  assign _T_2923 = releaseRejected ? 2'h0 : _T_2922; // @[DCache.scala 726:52]
  assign _GEN_350 = {{8'd0}, _T_2923}; // @[DCache.scala 726:47]
  assign releaseDataBeat = _T_2919 + _GEN_350; // @[DCache.scala 726:47]
  assign _T_2928 = s2_valid_flush_line | s2_flush_valid; // @[DCache.scala 739:34]
  assign _T_2929 = _T_2928 | io_cpu_s2_nack; // @[DCache.scala 739:52]
  assign _T_2931 = _T_2929 | reset; // @[DCache.scala 739:13]
  assign discard_line = s2_valid_flush_line & s2_req_size[1]; // @[DCache.scala 740:46]
  assign _T_2938 = s2_victim_dirty & ~discard_line; // @[DCache.scala 741:44]
  assign _T_2939 = _T_2938 ? 3'h1 : 3'h6; // @[DCache.scala 741:27]
  assign _T_2941 = {s2_victim_tag,s2_req_addr[11:6]}; // @[Cat.scala 29:58]
  assign res_2_address = {_T_2941, 6'h0}; // @[DCache.scala 742:96]
  assign _GEN_243 = s2_want_victimize ? _T_2939 : release_state; // @[DCache.scala 738:25]
  assign _T_2944 = releaseDone ? 3'h7 : 3'h3; // @[DCache.scala 753:29]
  assign _T_2946 = releaseDone ? 3'h0 : 3'h5; // @[DCache.scala 757:29]
  assign _GEN_254 = _T_2943 ? s2_report_param : 3'h5; // @[DCache.scala 750:45]
  assign _GEN_260 = _T_2943 ? _T_2944 : _T_2946; // @[DCache.scala 750:45]
  assign _GEN_262 = s2_prb_ack_data ? 3'h2 : _GEN_260; // @[DCache.scala 748:36]
  assign _GEN_265 = s2_prb_ack_data ? 3'h5 : _GEN_254; // @[DCache.scala 748:36]
  assign _GEN_272 = s2_meta_error ? 3'h4 : _GEN_262; // @[DCache.scala 746:28]
  assign _GEN_275 = s2_meta_error ? 3'h5 : _GEN_265; // @[DCache.scala 746:28]
  assign _GEN_283 = s2_probe ? _GEN_272 : _GEN_243; // @[DCache.scala 744:21]
  assign _GEN_286 = s2_probe ? _GEN_275 : 3'h5; // @[DCache.scala 744:21]
  assign _T_2947 = release_state == 3'h4; // @[DCache.scala 761:25]
  assign _T_2950 = {io_cpu_req_bits_addr[39:32],probe_bits_address}; // @[Cat.scala 29:58]
  assign _GEN_293 = metaArb_io_in_6_ready ? 3'h0 : _GEN_283; // @[DCache.scala 765:37]
  assign _GEN_294 = metaArb_io_in_6_ready | _T_17; // @[DCache.scala 765:37]
  assign _GEN_298 = _T_2947 ? _GEN_293 : _GEN_283; // @[DCache.scala 761:44]
  assign _GEN_300 = releaseDone ? 3'h0 : _GEN_298; // @[DCache.scala 772:26]
  assign _GEN_302 = _T_2951 ? _GEN_300 : _GEN_298; // @[DCache.scala 770:47]
  assign _GEN_306 = _T_2952 ? s2_report_param : _GEN_286; // @[DCache.scala 774:48]
  assign _GEN_315 = _T_2953 ? s2_report_param : _GEN_306; // @[DCache.scala 779:48]
  assign _T_2978 = _T_2898 & c_first; // @[DCache.scala 792:29]
  assign _GEN_323 = _T_2978 | _GEN_230; // @[DCache.scala 792:41]
  assign newCoh_state = _T_2956 ? voluntaryNewCoh_state : probeNewCoh_state; // @[DCache.scala 783:81]
  assign _T_2980 = releaseDataBeat < 10'h8; // @[DCache.scala 803:60]
  assign _T_2983 = {probe_bits_address[11:6], 6'h0}; // @[DCache.scala 806:55]
  assign _T_2985 = {releaseDataBeat[2:0], 3'h0}; // @[DCache.scala 806:117]
  assign _GEN_352 = {{6'd0}, _T_2985}; // @[DCache.scala 806:72]
  assign _T_2990 = release_state == 3'h7; // @[package.scala 15:47]
  assign _T_2999 = metaArb_io_in_4_ready & metaArb_io_in_4_valid; // @[Decoupled.scala 40:37]
  assign _T_3006 = s1_valid | s2_valid; // @[DCache.scala 829:57]
  assign _T_3007 = _T_3006 | cached_grant_wait; // @[DCache.scala 829:94]
  assign _T_3009 = _T_3007 | _T_661; // @[DCache.scala 829:115]
  assign _T_3012 = tlb_io_req_valid; // @[DCache.scala 831:40]
  assign _T_3027 = ~s2_valid_hit_pre_data_ecc_and_waw | reset; // @[DCache.scala 851:11]
  assign _T_3035 = s2_req_addr[2] ? s2_data_corrected[63:32] : s2_data_corrected[31:0]; // @[AMOALU.scala 39:24]
  assign _T_3038 = s2_req_size == 2'h2; // @[AMOALU.scala 42:26]
  assign _T_3041 = s2_req_signed & _T_3035[31]; // @[AMOALU.scala 42:76]
  assign _T_3043 = _T_3041 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _T_3045 = _T_3038 ? _T_3043 : s2_data_corrected[63:32]; // @[AMOALU.scala 42:20]
  assign _T_3046 = {_T_3045,_T_3035}; // @[Cat.scala 29:58]
  assign _T_3050 = s2_req_addr[1] ? _T_3046[31:16] : _T_3046[15:0]; // @[AMOALU.scala 39:24]
  assign _T_3053 = s2_req_size == 2'h1; // @[AMOALU.scala 42:26]
  assign _T_3056 = s2_req_signed & _T_3050[15]; // @[AMOALU.scala 42:76]
  assign _T_3058 = _T_3056 ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  assign _T_3060 = _T_3053 ? _T_3058 : _T_3046[63:16]; // @[AMOALU.scala 42:20]
  assign _T_3061 = {_T_3060,_T_3050}; // @[Cat.scala 29:58]
  assign _T_3065 = s2_req_addr[0] ? _T_3061[15:8] : _T_3061[7:0]; // @[AMOALU.scala 39:24]
  assign _T_3067 = _T_421 ? 8'h0 : _T_3065; // @[AMOALU.scala 41:23]
  assign _T_3068 = s2_req_size == 2'h0; // @[AMOALU.scala 42:26]
  assign _T_3069 = _T_3068 | _T_421; // @[AMOALU.scala 42:38]
  assign _T_3071 = s2_req_signed & _T_3067[7]; // @[AMOALU.scala 42:76]
  assign _T_3073 = _T_3071 ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  assign _T_3075 = _T_3069 ? _T_3073 : _T_3061[63:8]; // @[AMOALU.scala 42:20]
  assign _T_3076 = {_T_3075,_T_3067}; // @[Cat.scala 29:58]
  assign _GEN_353 = {{63'd0}, s2_sc_fail}; // @[DCache.scala 873:41]
  assign _GEN_341 = _T_3097 | resetting; // @[DCache.scala 908:27]
  assign flushCounterNext = flushCounter + 8'h1; // @[DCache.scala 910:39]
  assign flushDone = flushCounterNext[8:6] == 3'h4; // @[DCache.scala 911:57]
  assign _T_3103 = metaArb_io_in_5_ready & metaArb_io_in_5_valid; // @[Decoupled.scala 40:37]
  assign _T_3105 = _T_3103 & ~s1_flush_valid; // @[DCache.scala 915:45]
  assign _T_3107 = _T_3105 & ~s2_flush_valid_pre_tag_ecc; // @[DCache.scala 915:64]
  assign _T_3109 = _T_3107 & _T_78; // @[DCache.scala 915:95]
  assign _T_3116 = {metaArb_io_in_5_bits_idx, 6'h0}; // @[DCache.scala 919:98]
  assign _GEN_343 = resetting ? flushCounterNext : {{1'd0}, flushCounter}; // @[DCache.scala 952:20]
  assign _T_3180 = _T_3178 - 9'h1; // @[Edges.scala 231:28]
  assign _T_3181 = _T_3178 == 9'h0; // @[Edges.scala 232:25]
  assign _T_3182 = _T_3178 == 9'h1; // @[Edges.scala 233:25]
  assign _T_3184 = _T_3182 | _T_2910; // @[Edges.scala 233:37]
  assign auto_out_a_valid = s2_valid_uncached_pending | _T_2600; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_opcode = s2_uncached ? _T_2695_opcode : 3'h6; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_param = s2_uncached ? _T_2695_param : _T_2625_param; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_size = s2_uncached ? _T_2695_size : 4'h6; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_source = s2_uncached ? _T_2695_source : 1'h0; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_address = s2_uncached ? _T_2695_address : acquire_address[31:0]; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_mask = s2_uncached ? _T_2695_mask : 8'hff; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_data = s2_uncached ? _T_2695_data : 64'h0; // @[LazyModule.scala 305:12]
  assign auto_out_b_ready = metaArb_io_in_6_ready & ~_T_2892; // @[LazyModule.scala 305:12]
  assign auto_out_c_valid = _T_2952 | _GEN_301; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_opcode = _T_2956 ? 3'h7 : _GEN_314; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_param = _T_2956 ? s2_shrink_param : _GEN_315; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_size = _T_2956 ? 4'h6 : probe_bits_size; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_source = probe_bits_source; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_address = probe_bits_address; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_data = {_T_636,_T_633}; // @[LazyModule.scala 305:12]
  assign auto_out_d_ready = _T_2878 ? 1'h0 : _GEN_232; // @[LazyModule.scala 305:12]
  assign auto_out_e_valid = _T_2792 ? 1'h0 : _T_2779; // @[LazyModule.scala 305:12]
  assign auto_out_e_bits_sink = auto_out_d_bits_sink; // @[LazyModule.scala 305:12]
  assign io_cpu_req_ready = _T_2878 ? _GEN_233 : _GEN_31; // @[DCache.scala 203:20 DCache.scala 218:64 DCache.scala 226:53 DCache.scala 234:98 DCache.scala 699:26]
  assign io_cpu_s2_nack = _T_820 & ~s2_valid_hit_pre_data_ecc_and_waw; // @[DCache.scala 396:18]
  assign io_cpu_resp_valid = s2_valid_hit_pre_data_ecc_and_waw | doUncachedResp; // @[DCache.scala 848:21]
  assign io_cpu_resp_bits_tag = s2_req_tag; // @[DCache.scala 819:20]
  assign io_cpu_resp_bits_size = s2_req_size; // @[DCache.scala 819:20]
  assign io_cpu_resp_bits_data = _T_3076 | _GEN_353; // @[DCache.scala 819:20 DCache.scala 873:25]
  assign io_cpu_resp_bits_replay = doUncachedResp; // @[DCache.scala 821:27 DCache.scala 852:29]
  assign io_cpu_resp_bits_has_data = _T_400 | _T_439; // @[DCache.scala 820:29]
  assign io_cpu_resp_bits_data_word_bypass = {_T_3045,_T_3035}; // @[DCache.scala 874:37]
  assign io_cpu_replay_next = _T_2761 & grantIsUncachedData; // @[DCache.scala 849:22]
  assign io_cpu_s2_xcpt_ma_ld = _T_3014 & s2_tlb_xcpt_ma_ld; // @[DCache.scala 832:18]
  assign io_cpu_s2_xcpt_ma_st = _T_3014 & s2_tlb_xcpt_ma_st; // @[DCache.scala 832:18]
  assign io_cpu_s2_xcpt_pf_ld = _T_3014 & s2_tlb_xcpt_pf_ld; // @[DCache.scala 832:18]
  assign io_cpu_s2_xcpt_pf_st = _T_3014 & s2_tlb_xcpt_pf_st; // @[DCache.scala 832:18]
  assign io_cpu_s2_xcpt_ae_ld = _T_3014 & s2_tlb_xcpt_ae_ld; // @[DCache.scala 832:18]
  assign io_cpu_s2_xcpt_ae_st = _T_3014 & s2_tlb_xcpt_ae_st; // @[DCache.scala 832:18]
  assign io_cpu_ordered = ~_T_3009; // @[DCache.scala 829:18]
  assign io_cpu_perf_release = _T_3184 & _T_2898; // @[DCache.scala 978:23]
  assign io_cpu_perf_grant = auto_out_d_valid & d_last; // @[DCache.scala 979:21]
  assign io_ptw_req_valid = tlb_io_ptw_req_valid; // @[DCache.scala 230:10]
  assign io_ptw_req_bits_bits_addr = tlb_io_ptw_req_bits_bits_addr; // @[DCache.scala 230:10]
  assign tlb_clock = gated_clock;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = s1_valid_masked & s1_cmd_uses_tlb; // @[DCache.scala 232:20]
  assign tlb_io_req_bits_vaddr = s1_tlb_req_vaddr; // @[DCache.scala 233:19]
  assign tlb_io_req_bits_passthrough = s1_tlb_req_passthrough; // @[DCache.scala 233:19]
  assign tlb_io_req_bits_size = s1_tlb_req_size; // @[DCache.scala 233:19]
  assign tlb_io_req_bits_cmd = s1_tlb_req_cmd; // @[DCache.scala 233:19]
  assign tlb_io_sfence_valid = s1_valid_masked & s1_sfence; // @[DCache.scala 237:23]
  assign tlb_io_sfence_bits_rs1 = s1_req_size[0]; // @[DCache.scala 238:26]
  assign tlb_io_sfence_bits_rs2 = s1_req_size[1]; // @[DCache.scala 239:26]
  assign tlb_io_sfence_bits_addr = s1_req_addr[38:0]; // @[DCache.scala 241:27]
  assign tlb_io_ptw_req_ready = io_ptw_req_ready; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_ae = io_ptw_resp_bits_ae; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_level = io_ptw_resp_bits_level; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_homogeneous = io_ptw_resp_bits_homogeneous; // @[DCache.scala 230:10]
  assign tlb_io_ptw_ptbr_mode = io_ptw_ptbr_mode; // @[DCache.scala 230:10]
  assign tlb_io_ptw_status_debug = io_ptw_status_debug; // @[DCache.scala 230:10]
  assign tlb_io_ptw_status_dprv = io_ptw_status_dprv; // @[DCache.scala 230:10]
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_status_sum = io_ptw_status_sum; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask; // @[DCache.scala 230:10]
  assign pma_checker_clock = gated_clock;
  assign pma_checker_reset = reset;
  assign pma_checker_io_req_valid = 1'h0;
  assign pma_checker_io_req_bits_vaddr = 40'h0;
  assign pma_checker_io_req_bits_passthrough = 1'h1; // @[DCache.scala 247:39]
  assign pma_checker_io_req_bits_size = s1_req_size; // @[DCache.scala 248:27]
  assign pma_checker_io_req_bits_cmd = s1_req_cmd; // @[DCache.scala 248:27]
  assign pma_checker_io_sfence_valid = 1'h0;
  assign pma_checker_io_sfence_bits_rs1 = 1'h0;
  assign pma_checker_io_sfence_bits_rs2 = 1'h0;
  assign pma_checker_io_sfence_bits_addr = 39'h0;
  assign pma_checker_io_ptw_req_ready = 1'h0;
  assign pma_checker_io_ptw_resp_valid = 1'h0;
  assign pma_checker_io_ptw_resp_bits_ae = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_ppn = 54'h0;
  assign pma_checker_io_ptw_resp_bits_pte_d = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_a = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_g = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_u = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_x = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_w = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_r = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_v = 1'h0;
  assign pma_checker_io_ptw_resp_bits_level = 2'h0;
  assign pma_checker_io_ptw_resp_bits_homogeneous = 1'h0;
  assign pma_checker_io_ptw_ptbr_mode = 4'h0;
  assign pma_checker_io_ptw_status_debug = 1'h0;
  assign pma_checker_io_ptw_status_dprv = 2'h0;
  assign pma_checker_io_ptw_status_mxr = 1'h0;
  assign pma_checker_io_ptw_status_sum = 1'h0;
  assign pma_checker_io_ptw_pmp_0_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_0_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_0_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_0_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_0_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_0_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_0_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_1_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_1_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_1_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_1_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_1_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_1_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_1_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_2_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_2_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_2_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_2_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_2_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_2_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_2_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_3_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_3_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_3_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_3_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_3_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_3_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_3_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_4_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_4_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_4_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_4_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_4_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_4_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_4_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_5_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_5_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_5_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_5_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_5_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_5_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_5_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_6_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_6_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_6_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_6_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_6_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_6_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_6_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_7_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_7_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_7_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_7_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_7_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_7_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_7_mask = 32'h0;
  assign MaxPeriodFibonacciLFSR_clock = gated_clock;
  assign MaxPeriodFibonacciLFSR_reset = reset;
  assign MaxPeriodFibonacciLFSR_io_increment = _T_2761 & _GEN_208; // @[PRNG.scala 85:23]
  assign metaArb_io_in_0_valid = resetting; // @[DCache.scala 947:26]
  assign metaArb_io_in_0_bits_addr = metaArb_io_in_5_bits_addr; // @[DCache.scala 948:25]
  assign metaArb_io_in_0_bits_idx = metaArb_io_in_5_bits_idx; // @[DCache.scala 948:25]
  assign metaArb_io_in_0_bits_data = {2'h0,s2_req_addr[31:12]}; // @[DCache.scala 948:25 DCache.scala 951:30]
  assign metaArb_io_in_1_valid = s2_meta_error & _T_832; // @[DCache.scala 401:26]
  assign metaArb_io_in_1_bits_addr = {io_cpu_req_bits_addr[39:12],_T_848}; // @[DCache.scala 405:30]
  assign metaArb_io_in_1_bits_idx = s2_probe ? probe_bits_address[11:6] : s2_vaddr[11:6]; // @[DCache.scala 404:29]
  assign metaArb_io_in_1_bits_data = {new_meta_coh_state,s2_meta_corrected_3_tag}; // @[DCache.scala 406:30]
  assign metaArb_io_in_2_valid = s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta; // @[DCache.scala 413:26]
  assign metaArb_io_in_2_bits_addr = {io_cpu_req_bits_addr[39:12],s2_vaddr[11:0]}; // @[DCache.scala 417:30]
  assign metaArb_io_in_2_bits_idx = s2_vaddr[11:6]; // @[DCache.scala 416:29]
  assign metaArb_io_in_2_bits_way_en = s2_hit_valid ? s2_hit_way : _T_673; // @[DCache.scala 415:32]
  assign metaArb_io_in_2_bits_data = {s2_grow_param,s2_req_addr[31:12]}; // @[DCache.scala 418:30]
  assign metaArb_io_in_3_valid = _T_2798 & ~auto_out_d_bits_denied; // @[DCache.scala 684:26]
  assign metaArb_io_in_3_bits_addr = {io_cpu_req_bits_addr[39:12],s2_vaddr[11:0]}; // @[DCache.scala 688:30]
  assign metaArb_io_in_3_bits_idx = s2_vaddr[11:6]; // @[DCache.scala 687:29]
  assign metaArb_io_in_3_bits_way_en = s2_hit_valid ? s2_hit_way : _T_673; // @[DCache.scala 686:32]
  assign metaArb_io_in_3_bits_data = {_T_2873,s2_req_addr[31:12]}; // @[DCache.scala 689:30]
  assign metaArb_io_in_4_valid = _T_2955 | _T_2990; // @[DCache.scala 810:26]
  assign metaArb_io_in_4_bits_addr = {io_cpu_req_bits_addr[39:12],probe_bits_address[11:0]}; // @[DCache.scala 814:30]
  assign metaArb_io_in_4_bits_idx = probe_bits_address[11:6]; // @[DCache.scala 813:29]
  assign metaArb_io_in_4_bits_way_en = _T_2956 ? s2_victim_way : s2_probe_way; // @[DCache.scala 812:32]
  assign metaArb_io_in_4_bits_data = {newCoh_state,probe_bits_address[31:12]}; // @[DCache.scala 815:30]
  assign metaArb_io_in_5_valid = 1'h0; // @[DCache.scala 916:26]
  assign metaArb_io_in_5_bits_addr = {io_cpu_req_bits_addr[39:12],_T_3116}; // @[DCache.scala 919:30]
  assign metaArb_io_in_5_bits_idx = flushCounter[5:0]; // @[DCache.scala 918:29]
  assign metaArb_io_in_6_valid = _T_2947 | _T_2889; // @[DCache.scala 712:26 DCache.scala 762:30]
  assign metaArb_io_in_6_bits_addr = _T_2947 ? _T_2950 : _T_2897; // @[DCache.scala 716:30 DCache.scala 764:34]
  assign metaArb_io_in_6_bits_idx = _T_2947 ? probe_bits_address[11:6] : auto_out_b_bits_address[11:6]; // @[DCache.scala 715:29 DCache.scala 763:33]
  assign metaArb_io_in_6_bits_way_en = metaArb_io_in_4_bits_way_en; // @[DCache.scala 717:32]
  assign metaArb_io_in_6_bits_data = metaArb_io_in_4_bits_data; // @[DCache.scala 718:30]
  assign metaArb_io_in_7_valid = io_cpu_req_valid; // @[DCache.scala 220:26]
  assign metaArb_io_in_7_bits_addr = io_cpu_req_bits_addr; // @[DCache.scala 223:30]
  assign metaArb_io_in_7_bits_idx = io_cpu_req_bits_addr[11:6]; // @[DCache.scala 222:29]
  assign metaArb_io_in_7_bits_way_en = metaArb_io_in_4_bits_way_en; // @[DCache.scala 224:32]
  assign metaArb_io_in_7_bits_data = metaArb_io_in_4_bits_data; // @[DCache.scala 225:30]
  assign data_clock = gated_clock;
  assign data_io_req_valid = dataArb_io_out_valid; // @[DCache.scala 133:15]
  assign data_io_req_bits_addr = dataArb_io_out_bits_addr; // @[DCache.scala 133:15]
  assign data_io_req_bits_write = dataArb_io_out_bits_write; // @[DCache.scala 133:15]
  assign data_io_req_bits_wdata = dataArb_io_out_bits_wdata; // @[DCache.scala 133:15]
  assign data_io_req_bits_eccMask = dataArb_io_out_bits_eccMask; // @[DCache.scala 133:15]
  assign data_io_req_bits_way_en = dataArb_io_out_bits_way_en; // @[DCache.scala 133:15]
  assign dataArb_io_in_0_valid = pstore_drain_structural | _T_1048; // @[DCache.scala 498:26]
  assign dataArb_io_in_0_bits_addr = _T_1132[11:0]; // @[DCache.scala 500:30]
  assign dataArb_io_in_0_bits_write = pstore_drain_structural | _T_1048; // @[DCache.scala 499:31]
  assign dataArb_io_in_0_bits_wdata = {_T_1148,_T_1145}; // @[DCache.scala 502:31]
  assign dataArb_io_in_0_bits_eccMask = {_T_1174,_T_1171}; // @[DCache.scala 504:33]
  assign dataArb_io_in_0_bits_way_en = pstore2_valid ? pstore2_way : pstore1_way; // @[DCache.scala 501:32]
  assign dataArb_io_in_1_valid = _T_2878 ? _GEN_234 : _T_2790; // @[DCache.scala 664:26 DCache.scala 700:32]
  assign dataArb_io_in_1_bits_addr = _T_2795[11:0]; // @[DCache.scala 671:32]
  assign dataArb_io_in_1_bits_write = _T_2878 ? _GEN_235 : 1'h1; // @[DCache.scala 670:33 DCache.scala 701:37]
  assign dataArb_io_in_1_bits_wdata = {_T_335,_T_332}; // @[DCache.scala 132:43 DCache.scala 673:33]
  assign dataArb_io_in_1_bits_eccMask = 8'hff; // @[DCache.scala 675:35]
  assign dataArb_io_in_1_bits_way_en = s2_hit_valid ? s2_hit_way : _T_673; // @[DCache.scala 672:34]
  assign dataArb_io_in_2_valid = inWriteback & _T_2980; // @[DCache.scala 803:26]
  assign dataArb_io_in_2_bits_addr = _T_2983 | _GEN_352; // @[DCache.scala 804:25 DCache.scala 806:30]
  assign dataArb_io_in_2_bits_wdata = dataArb_io_in_1_bits_wdata; // @[DCache.scala 132:43 DCache.scala 804:25]
  assign dataArb_io_in_2_bits_eccMask = dataArb_io_in_1_bits_eccMask; // @[DCache.scala 804:25]
  assign dataArb_io_in_3_valid = io_cpu_req_valid & res; // @[DCache.scala 212:26]
  assign dataArb_io_in_3_bits_addr = io_cpu_req_bits_addr[11:0]; // @[DCache.scala 213:25 DCache.scala 215:30]
  assign dataArb_io_in_3_bits_wdata = dataArb_io_in_1_bits_wdata; // @[DCache.scala 132:43 DCache.scala 213:25]
  assign dataArb_io_in_3_bits_eccMask = dataArb_io_in_1_bits_eccMask; // @[DCache.scala 213:25]
  assign amoalu_io_mask = pstore1_mask; // @[DCache.scala 882:22]
  assign amoalu_io_cmd = pstore1_cmd; // @[DCache.scala 883:21]
  assign amoalu_io_lhs = {_T_636,_T_633}; // @[DCache.scala 884:21]
  assign amoalu_io_rhs = pstore1_data; // @[DCache.scala 885:21]
  assign _GEN_356 = _T_2761 & grantIsCached; // @[DCache.scala 620:13]
  assign _GEN_359 = _T_2761 & ~grantIsCached; // @[DCache.scala 630:17]
  assign _GEN_360 = _GEN_359 & grantIsUncached; // @[DCache.scala 630:17]
  assign _GEN_361 = _GEN_360 & _T_2766; // @[DCache.scala 630:17]
  assign _GEN_369 = _GEN_359 & ~grantIsUncached; // @[DCache.scala 651:13]
  assign _GEN_370 = _GEN_369 & grantIsVoluntary; // @[DCache.scala 651:13]
  assign DCache_cov_read_addr = DCache_state;
  assign DCache_cov_read_data = DCache_cov[DCache_cov_read_addr]; // @[Coverage map for DCache]
  assign DCache_cov_write_data = 1'h1;
  assign DCache_cov_write_addr = DCache_state;
  assign DCache_cov_write_mask = 1'h1;
  assign DCache_cov_write_en = 1'h1;
  assign mux_cond_0 = s1_req_addr[0];
  assign mux_cond_1 = s2_req_addr[0];
  assign mux_cond_2 = s2_req_addr[1];
  assign mux_cond_3 = s1_req_addr[1];
  assign mux_cond_4 = s1_req_addr[2];
  assign mux_cond_5 = s2_req_addr[2];
  assign pstore1_held_shl = {pstore1_held, 9'h0};
  assign pstore1_held_pad = {10'h0,pstore1_held_shl};
  assign pstore2_valid_shl = {pstore2_valid, 5'h0};
  assign pstore2_valid_pad = {14'h0,pstore2_valid_shl};
  assign s2_valid_shl = {s2_valid, 2'h0};
  assign s2_valid_pad = {17'h0,s2_valid_shl};
  assign release_state_shl = {release_state, 15'h0};
  assign release_state_pad = {2'h0,release_state_shl};
  assign s2_probe_shl = {s2_probe, 7'h0};
  assign s2_probe_pad = {12'h0,s2_probe_shl};
  assign s2_flush_valid_pre_tag_ecc_shl = s2_flush_valid_pre_tag_ecc;
  assign s2_flush_valid_pre_tag_ecc_pad = {19'h0,s2_flush_valid_pre_tag_ecc_shl};
  assign _T_679_state_shl = {_T_679_state, 9'h0};
  assign _T_679_state_pad = {9'h0,_T_679_state_shl};
  assign uncachedInFlight_0_shl = {uncachedInFlight_0, 1'h0};
  assign uncachedInFlight_0_pad = {18'h0,uncachedInFlight_0_shl};
  assign s2_release_data_valid_shl = {s2_release_data_valid, 14'h0};
  assign s2_release_data_valid_pad = {5'h0,s2_release_data_valid_shl};
  assign probe_bits_param_shl = {probe_bits_param, 6'h0};
  assign probe_bits_param_pad = {12'h0,probe_bits_param_shl};
  assign s2_pma_cacheable_shl = {s2_pma_cacheable, 14'h0};
  assign s2_pma_cacheable_pad = {5'h0,s2_pma_cacheable_shl};
  assign s2_hit_state_state_shl = {s2_hit_state_state, 12'h0};
  assign s2_hit_state_state_pad = {6'h0,s2_hit_state_state_shl};
  assign s2_req_size_shl = s2_req_size;
  assign s2_req_size_pad = {18'h0,s2_req_size_shl};
  assign s1_did_read_shl = s1_did_read;
  assign s1_did_read_pad = {19'h0,s1_did_read_shl};
  assign grantInProgress_shl = {grantInProgress, 11'h0};
  assign grantInProgress_pad = {8'h0,grantInProgress_shl};
  assign _T_1016_shl = {_T_1016, 11'h0};
  assign _T_1016_pad = {8'h0,_T_1016_shl};
  assign s2_not_nacked_in_s1_shl = {s2_not_nacked_in_s1, 12'h0};
  assign s2_not_nacked_in_s1_pad = {7'h0,s2_not_nacked_in_s1_shl};
  assign blockUncachedGrant_shl = {blockUncachedGrant, 19'h0};
  assign blockUncachedGrant_pad = blockUncachedGrant_shl;
  assign _T_672_shl = {_T_672, 15'h0};
  assign _T_672_pad = {3'h0,_T_672_shl};
  assign s2_hit_way_shl = {s2_hit_way, 3'h0};
  assign s2_hit_way_pad = {13'h0,s2_hit_way_shl};
  assign cached_grant_wait_shl = {cached_grant_wait, 19'h0};
  assign cached_grant_wait_pad = cached_grant_wait_shl;
  assign s2_req_signed_shl = {s2_req_signed, 11'h0};
  assign s2_req_signed_pad = {8'h0,s2_req_signed_shl};
  assign release_ack_wait_shl = {release_ack_wait, 16'h0};
  assign release_ack_wait_pad = {3'h0,release_ack_wait_shl};
  assign s2_probe_state_state_shl = {s2_probe_state_state, 2'h0};
  assign s2_probe_state_state_pad = {16'h0,s2_probe_state_state_shl};
  assign s1_probe_shl = {s1_probe, 2'h0};
  assign s1_probe_pad = {17'h0,s1_probe_shl};
  assign s1_valid_shl = {s1_valid, 1'h0};
  assign s1_valid_pad = {18'h0,s1_valid_shl};
  assign s1_req_size_shl = {s1_req_size, 5'h0};
  assign s1_req_size_pad = {13'h0,s1_req_size_shl};
  assign pstore1_rmw_shl = {pstore1_rmw, 15'h0};
  assign pstore1_rmw_pad = {4'h0,pstore1_rmw_shl};
  assign s1_flush_valid_shl = {s1_flush_valid, 11'h0};
  assign s1_flush_valid_pad = {8'h0,s1_flush_valid_shl};
  assign resetting_shl = resetting;
  assign resetting_pad = {19'h0,resetting_shl};
  assign s2_probe_way_shl = {s2_probe_way, 12'h0};
  assign s2_probe_way_pad = {4'h0,s2_probe_way_shl};
  assign mux_cond_0_shl = {mux_cond_0, 9'h0};
  assign mux_cond_0_pad = {10'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 2'h0};
  assign mux_cond_1_pad = {17'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 7'h0};
  assign mux_cond_2_pad = {12'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 15'h0};
  assign mux_cond_3_pad = {4'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 5'h0};
  assign mux_cond_4_pad = {14'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 19'h0};
  assign mux_cond_5_pad = mux_cond_5_shl;
  assign DCache_xor15 = pstore1_held_pad ^ pstore2_valid_pad;
  assign DCache_xor16 = s2_valid_pad ^ release_state_pad;
  assign DCache_xor7 = DCache_xor15 ^ DCache_xor16;
  assign DCache_xor17 = s2_probe_pad ^ s2_flush_valid_pre_tag_ecc_pad;
  assign DCache_xor38 = uncachedInFlight_0_pad ^ s2_release_data_valid_pad;
  assign DCache_xor18 = _T_679_state_pad ^ DCache_xor38;
  assign DCache_xor8 = DCache_xor17 ^ DCache_xor18;
  assign DCache_xor3 = DCache_xor7 ^ DCache_xor8;
  assign DCache_xor19 = probe_bits_param_pad ^ s2_pma_cacheable_pad;
  assign DCache_xor20 = s2_hit_state_state_pad ^ s2_req_size_pad;
  assign DCache_xor9 = DCache_xor19 ^ DCache_xor20;
  assign DCache_xor21 = s1_did_read_pad ^ grantInProgress_pad;
  assign DCache_xor46 = s2_not_nacked_in_s1_pad ^ blockUncachedGrant_pad;
  assign DCache_xor22 = _T_1016_pad ^ DCache_xor46;
  assign DCache_xor10 = DCache_xor21 ^ DCache_xor22;
  assign DCache_xor4 = DCache_xor9 ^ DCache_xor10;
  assign DCache_xor1 = DCache_xor3 ^ DCache_xor4;
  assign DCache_xor23 = _T_672_pad ^ s2_hit_way_pad;
  assign DCache_xor24 = cached_grant_wait_pad ^ s2_req_signed_pad;
  assign DCache_xor11 = DCache_xor23 ^ DCache_xor24;
  assign DCache_xor25 = release_ack_wait_pad ^ s2_probe_state_state_pad;
  assign DCache_xor54 = s1_valid_pad ^ s1_req_size_pad;
  assign DCache_xor26 = s1_probe_pad ^ DCache_xor54;
  assign DCache_xor12 = DCache_xor25 ^ DCache_xor26;
  assign DCache_xor5 = DCache_xor11 ^ DCache_xor12;
  assign DCache_xor27 = pstore1_rmw_pad ^ s1_flush_valid_pad;
  assign DCache_xor58 = s2_probe_way_pad ^ mux_cond_0_pad;
  assign DCache_xor28 = resetting_pad ^ DCache_xor58;
  assign DCache_xor13 = DCache_xor27 ^ DCache_xor28;
  assign DCache_xor29 = mux_cond_1_pad ^ mux_cond_2_pad;
  assign DCache_xor62 = mux_cond_4_pad ^ mux_cond_5_pad;
  assign DCache_xor30 = mux_cond_3_pad ^ DCache_xor62;
  assign DCache_xor14 = DCache_xor29 ^ DCache_xor30;
  assign DCache_xor6 = DCache_xor13 ^ DCache_xor14;
  assign DCache_xor2 = DCache_xor5 ^ DCache_xor6;
  assign DCache_xor0 = DCache_xor1 ^ DCache_xor2;
  assign amoalu_sum = DCache_covSum + amoalu_io_covSum;
  assign MaxPeriodFibonacciLFSR_sum = amoalu_sum + MaxPeriodFibonacciLFSR_io_covSum;
  assign pma_checker_sum = MaxPeriodFibonacciLFSR_sum + pma_checker_io_covSum;
  assign metaArb_sum = pma_checker_sum + metaArb_io_covSum;
  assign dataArb_sum = metaArb_sum + dataArb_io_covSum;
  assign tlb_sum = dataArb_sum + tlb_io_covSum;
  assign data_sum = tlb_sum + data_io_covSum;
  assign io_covSum = data_sum;
  assign stopEn0 = ~_T_165;
  assign stopEn1 = ~_T_370;
  assign stopEn2 = ~_T_165;
  assign stopEn3 = ~_T_1034;
  assign stopEn4 = _GEN_356 & ~_T_2763;
  assign stopEn5 = _GEN_361 & ~_T_2768;
  assign stopEn6 = _GEN_370 & ~_T_2775;
  assign stopEn7 = ~_T_2787;
  assign stopEn8 = s2_want_victimize & ~_T_2931;
  assign stopEn9 = doUncachedResp & ~_T_3027;
  assign tlb_metaAssert_wire = tlb_metaAssert;
  assign amoalu_metaAssert_wire = amoalu_metaAssert;
  assign dataArb_metaAssert_wire = dataArb_metaAssert;
  assign metaArb_metaAssert_wire = metaArb_metaAssert;
  assign data_metaAssert_wire = data_metaAssert;
  assign MaxPeriodFibonacciLFSR_metaAssert_wire = MaxPeriodFibonacciLFSR_metaAssert;
  assign pma_checker_metaAssert_wire = pma_checker_metaAssert;
  assign DCache_or7 = stopEn0 | stopEn1;
  assign DCache_or8 = stopEn2 | stopEn3;
  assign DCache_or3 = DCache_or7 | DCache_or8;
  assign DCache_or9 = stopEn4 | stopEn5;
  assign DCache_or10 = stopEn6 | stopEn7;
  assign DCache_or4 = DCache_or9 | DCache_or10;
  assign DCache_or1 = DCache_or3 | DCache_or4;
  assign DCache_or11 = stopEn8 | stopEn9;
  assign DCache_or12 = dataArb_metaAssert_wire | MaxPeriodFibonacciLFSR_metaAssert_wire;
  assign DCache_or5 = DCache_or11 | DCache_or12;
  assign DCache_or13 = tlb_metaAssert_wire | amoalu_metaAssert_wire;
  assign DCache_or30 = pma_checker_metaAssert_wire | metaArb_metaAssert_wire;
  assign DCache_or14 = data_metaAssert_wire | DCache_or30;
  assign DCache_or6 = DCache_or13 | DCache_or14;
  assign DCache_or2 = DCache_or5 | DCache_or6;
  assign DCache_or0 = DCache_or1 | DCache_or2;
  assign metaAssert = DCache_or0;
  assign MaxPeriodFibonacciLFSR_metaReset = metaReset | MaxPeriodFibonacciLFSR_halt;
  assign pma_checker_metaReset = metaReset | pma_checker_halt;
  assign tlb_metaReset = metaReset | tlb_halt;
  assign data_metaReset = metaReset | data_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_0[initvar] = _RAND_0[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tag_array_0_s1_meta_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tag_array_0_s1_meta_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_1[initvar] = _RAND_3[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  tag_array_1_s1_meta_en_pipe_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  tag_array_1_s1_meta_addr_pipe_0 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_2[initvar] = _RAND_6[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  tag_array_2_s1_meta_en_pipe_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tag_array_2_s1_meta_addr_pipe_0 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_3[initvar] = _RAND_9[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  tag_array_3_s1_meta_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  tag_array_3_s1_meta_addr_pipe_0 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  s1_valid = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  blockProbeAfterGrantCount = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  lrscCount = _RAND_14[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  s1_probe = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  s2_probe = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  release_state = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  release_ack_wait = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  release_ack_addr = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  grantInProgress = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  s2_valid = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  probe_bits_param = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  probe_bits_size = _RAND_23[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  probe_bits_source = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  probe_bits_address = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  s2_probe_state_state = _RAND_26[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_2906 = _RAND_27[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  s2_release_data_valid = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  s1_req_cmd = _RAND_29[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  s2_req_cmd = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  pstore1_held = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  pstore1_addr = _RAND_32[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{`RANDOM}};
  s1_req_addr = _RAND_33[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  pstore1_mask = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  s1_req_size = _RAND_35[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  pstore2_valid = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  pstore2_addr = _RAND_37[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  mask = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  s2_not_nacked_in_s1 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  s2_hit_state_state = _RAND_40[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  s1_req_tag = _RAND_41[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  s1_req_signed = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{`RANDOM}};
  s1_tlb_req_vaddr = _RAND_43[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  s1_tlb_req_passthrough = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  s1_tlb_req_size = _RAND_45[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  s1_tlb_req_cmd = _RAND_46[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  s1_flush_valid = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  cached_grant_wait = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  uncachedInFlight_0 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {2{`RANDOM}};
  uncachedReqs_0_addr = _RAND_50[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  uncachedReqs_0_tag = _RAND_51[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  uncachedReqs_0_size = _RAND_52[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  uncachedReqs_0_signed = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  s1_did_read = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  s2_hit_way = _RAND_55[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_672 = _RAND_56[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  s2_probe_way = _RAND_57[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  s2_req_addr = _RAND_58[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  s2_req_tag = _RAND_59[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  s2_req_size = _RAND_60[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  s2_req_signed = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  s2_tlb_xcpt_pf_ld = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  s2_tlb_xcpt_pf_st = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  s2_tlb_xcpt_ae_ld = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  s2_tlb_xcpt_ae_st = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  s2_tlb_xcpt_ma_ld = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  s2_tlb_xcpt_ma_st = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  s2_pma_cacheable = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {2{`RANDOM}};
  _T_393 = _RAND_69[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  s2_flush_valid_pre_tag_ecc = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_465 = _RAND_71[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  blockUncachedGrant = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_2713 = _RAND_73[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{`RANDOM}};
  s2_data = _RAND_74[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_677 = _RAND_75[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_679_state = _RAND_76[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {2{`RANDOM}};
  lrscAddr = _RAND_77[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  pstore1_cmd = _RAND_78[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {2{`RANDOM}};
  pstore1_data = _RAND_79[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  pstore1_way = _RAND_80[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  pstore1_rmw = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_1016 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  pstore2_way = _RAND_83[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_1072 = _RAND_84[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_1077 = _RAND_85[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_1082 = _RAND_86[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_1087 = _RAND_87[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_1092 = _RAND_88[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_1097 = _RAND_89[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_1102 = _RAND_90[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_1107 = _RAND_91[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  s1_release_data_valid = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_3014 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  doUncachedResp = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  resetting = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_3097 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  flushCounter = _RAND_97[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_3178 = _RAND_98[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  DCache_state = _RAND_99[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    DCache_cov[initvar] = _RAND_100[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  DCache_covSum = _RAND_101[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge gated_clock) begin
    if(tag_array_0__T_260_en & tag_array_0__T_260_mask) begin
      tag_array_0[tag_array_0__T_260_addr] <= tag_array_0__T_260_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      tag_array_0_s1_meta_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_0_s1_meta_en_pipe_0 <= metaArb_io_out_valid & ~metaArb_io_out_bits_write;
    end
    if (metaReset) begin
      tag_array_0_s1_meta_addr_pipe_0 <= 6'h0;
    end else if (metaArb_io_out_valid & ~metaArb_io_out_bits_write) begin
      tag_array_0_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if(tag_array_1__T_260_en & tag_array_1__T_260_mask) begin
      tag_array_1[tag_array_1__T_260_addr] <= tag_array_1__T_260_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      tag_array_1_s1_meta_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_1_s1_meta_en_pipe_0 <= metaArb_io_out_valid & ~metaArb_io_out_bits_write;
    end
    if (metaReset) begin
      tag_array_1_s1_meta_addr_pipe_0 <= 6'h0;
    end else if (metaArb_io_out_valid & ~metaArb_io_out_bits_write) begin
      tag_array_1_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if(tag_array_2__T_260_en & tag_array_2__T_260_mask) begin
      tag_array_2[tag_array_2__T_260_addr] <= tag_array_2__T_260_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      tag_array_2_s1_meta_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_2_s1_meta_en_pipe_0 <= metaArb_io_out_valid & ~metaArb_io_out_bits_write;
    end
    if (metaReset) begin
      tag_array_2_s1_meta_addr_pipe_0 <= 6'h0;
    end else if (metaArb_io_out_valid & ~metaArb_io_out_bits_write) begin
      tag_array_2_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if(tag_array_3__T_260_en & tag_array_3__T_260_mask) begin
      tag_array_3[tag_array_3__T_260_addr] <= tag_array_3__T_260_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      tag_array_3_s1_meta_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_3_s1_meta_en_pipe_0 <= metaArb_io_out_valid & ~metaArb_io_out_bits_write;
    end
    if (metaReset) begin
      tag_array_3_s1_meta_addr_pipe_0 <= 6'h0;
    end else if (metaArb_io_out_valid & ~metaArb_io_out_bits_write) begin
      tag_array_3_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if (metaReset) begin
      s1_valid <= 1'h0;
    end else if (reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= _T_16;
    end
    if (metaReset) begin
      blockProbeAfterGrantCount <= 3'h0;
    end else if (reset) begin
      blockProbeAfterGrantCount <= 3'h0;
    end else if (_T_2761) begin
      if (grantIsCached) begin
        if (d_last) begin
          blockProbeAfterGrantCount <= 3'h7;
        end else if (_T_2882) begin
          blockProbeAfterGrantCount <= _T_2749;
        end
      end else if (_T_2882) begin
        blockProbeAfterGrantCount <= _T_2749;
      end
    end else if (_T_2882) begin
      blockProbeAfterGrantCount <= _T_2749;
    end
    if (metaReset) begin
      lrscCount <= 7'h0;
    end else if (reset) begin
      lrscCount <= 7'h0;
    end else if (s1_probe) begin
      lrscCount <= 7'h0;
    end else if (_T_879) begin
      lrscCount <= 7'h3;
    end else if (_T_863) begin
      lrscCount <= _T_878;
    end else if (_T_871) begin
      if (s2_hit) begin
        lrscCount <= 7'h4f;
      end else begin
        lrscCount <= 7'h0;
      end
    end
    if (metaReset) begin
      s1_probe <= 1'h0;
    end else if (reset) begin
      s1_probe <= 1'h0;
    end else if (_T_2947) begin
      s1_probe <= _GEN_294;
    end else begin
      s1_probe <= _T_17;
    end
    if (metaReset) begin
      s2_probe <= 1'h0;
    end else if (reset) begin
      s2_probe <= 1'h0;
    end else begin
      s2_probe <= s1_probe;
    end
    if (metaReset) begin
      release_state <= 3'h0;
    end else if (reset) begin
      release_state <= 3'h0;
    end else if (_T_2999) begin
      release_state <= 3'h0;
    end else if (_T_2956) begin
      if (releaseDone) begin
        release_state <= 3'h6;
      end else if (_T_2953) begin
        if (releaseDone) begin
          release_state <= 3'h7;
        end else if (_T_2952) begin
          if (releaseDone) begin
            release_state <= 3'h7;
          end else if (_T_2951) begin
            if (releaseDone) begin
              release_state <= 3'h0;
            end else if (_T_2947) begin
              if (metaArb_io_in_6_ready) begin
                release_state <= 3'h0;
              end else if (s2_probe) begin
                if (s2_meta_error) begin
                  release_state <= 3'h4;
                end else if (s2_prb_ack_data) begin
                  release_state <= 3'h2;
                end else if (_T_2943) begin
                  if (releaseDone) begin
                    release_state <= 3'h7;
                  end else begin
                    release_state <= 3'h3;
                  end
                end else if (releaseDone) begin
                  release_state <= 3'h0;
                end else begin
                  release_state <= 3'h5;
                end
              end else if (s2_want_victimize) begin
                if (_T_2938) begin
                  release_state <= 3'h1;
                end else begin
                  release_state <= 3'h6;
                end
              end
            end else if (s2_probe) begin
              if (s2_meta_error) begin
                release_state <= 3'h4;
              end else if (s2_prb_ack_data) begin
                release_state <= 3'h2;
              end else if (_T_2943) begin
                if (releaseDone) begin
                  release_state <= 3'h7;
                end else begin
                  release_state <= 3'h3;
                end
              end else if (releaseDone) begin
                release_state <= 3'h0;
              end else begin
                release_state <= 3'h5;
              end
            end else if (s2_want_victimize) begin
              if (_T_2938) begin
                release_state <= 3'h1;
              end else begin
                release_state <= 3'h6;
              end
            end
          end else if (_T_2947) begin
            if (metaArb_io_in_6_ready) begin
              release_state <= 3'h0;
            end else if (s2_probe) begin
              if (s2_meta_error) begin
                release_state <= 3'h4;
              end else if (s2_prb_ack_data) begin
                release_state <= 3'h2;
              end else if (_T_2943) begin
                if (releaseDone) begin
                  release_state <= 3'h7;
                end else begin
                  release_state <= 3'h3;
                end
              end else if (releaseDone) begin
                release_state <= 3'h0;
              end else begin
                release_state <= 3'h5;
              end
            end else if (s2_want_victimize) begin
              if (_T_2938) begin
                release_state <= 3'h1;
              end else begin
                release_state <= 3'h6;
              end
            end
          end else if (s2_probe) begin
            if (s2_meta_error) begin
              release_state <= 3'h4;
            end else if (s2_prb_ack_data) begin
              release_state <= 3'h2;
            end else if (_T_2943) begin
              if (releaseDone) begin
                release_state <= 3'h7;
              end else begin
                release_state <= 3'h3;
              end
            end else if (releaseDone) begin
              release_state <= 3'h0;
            end else begin
              release_state <= 3'h5;
            end
          end else if (s2_want_victimize) begin
            if (_T_2938) begin
              release_state <= 3'h1;
            end else begin
              release_state <= 3'h6;
            end
          end
        end else if (_T_2951) begin
          if (releaseDone) begin
            release_state <= 3'h0;
          end else if (_T_2947) begin
            if (metaArb_io_in_6_ready) begin
              release_state <= 3'h0;
            end else begin
              release_state <= _GEN_283;
            end
          end else begin
            release_state <= _GEN_283;
          end
        end else if (_T_2947) begin
          if (metaArb_io_in_6_ready) begin
            release_state <= 3'h0;
          end else begin
            release_state <= _GEN_283;
          end
        end else begin
          release_state <= _GEN_283;
        end
      end else if (_T_2952) begin
        if (releaseDone) begin
          release_state <= 3'h7;
        end else if (_T_2951) begin
          if (releaseDone) begin
            release_state <= 3'h0;
          end else begin
            release_state <= _GEN_298;
          end
        end else begin
          release_state <= _GEN_298;
        end
      end else if (_T_2951) begin
        if (releaseDone) begin
          release_state <= 3'h0;
        end else begin
          release_state <= _GEN_298;
        end
      end else begin
        release_state <= _GEN_298;
      end
    end else if (_T_2953) begin
      if (releaseDone) begin
        release_state <= 3'h7;
      end else if (_T_2952) begin
        if (releaseDone) begin
          release_state <= 3'h7;
        end else begin
          release_state <= _GEN_302;
        end
      end else begin
        release_state <= _GEN_302;
      end
    end else if (_T_2952) begin
      if (releaseDone) begin
        release_state <= 3'h7;
      end else begin
        release_state <= _GEN_302;
      end
    end else begin
      release_state <= _GEN_302;
    end
    if (metaReset) begin
      release_ack_wait <= 1'h0;
    end else if (reset) begin
      release_ack_wait <= 1'h0;
    end else if (_T_2956) begin
      release_ack_wait <= _GEN_323;
    end else if (_T_2761) begin
      if (!(grantIsCached)) begin
        if (!(grantIsUncached)) begin
          if (grantIsVoluntary) begin
            release_ack_wait <= 1'h0;
          end
        end
      end
    end
    if (metaReset) begin
      release_ack_addr <= 32'h0;
    end else if (_T_2956) begin
      if (_T_2978) begin
        release_ack_addr <= probe_bits_address;
      end
    end
    if (metaReset) begin
      grantInProgress <= 1'h0;
    end else if (reset) begin
      grantInProgress <= 1'h0;
    end else if (_T_2761) begin
      if (grantIsCached) begin
        if (d_last) begin
          grantInProgress <= 1'h0;
        end else begin
          grantInProgress <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      s2_valid <= 1'h0;
    end else if (reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= _T_373;
    end
    if (metaReset) begin
      probe_bits_param <= 2'h0;
    end else if (s2_want_victimize) begin
      probe_bits_param <= 2'h0;
    end else if (_T_17) begin
      probe_bits_param <= auto_out_b_bits_param;
    end
    if (metaReset) begin
      probe_bits_size <= 4'h0;
    end else if (s2_want_victimize) begin
      probe_bits_size <= 4'h0;
    end else if (_T_17) begin
      probe_bits_size <= auto_out_b_bits_size;
    end
    if (metaReset) begin
      probe_bits_source <= 1'h0;
    end else if (s2_want_victimize) begin
      probe_bits_source <= 1'h0;
    end else if (_T_17) begin
      probe_bits_source <= auto_out_b_bits_source;
    end
    if (metaReset) begin
      probe_bits_address <= 32'h0;
    end else if (s2_want_victimize) begin
      probe_bits_address <= res_2_address;
    end else if (_T_17) begin
      probe_bits_address <= auto_out_b_bits_address;
    end
    if (metaReset) begin
      s2_probe_state_state <= 2'h0;
    end else if (s1_probe) begin
      s2_probe_state_state <= s1_meta_hit_state_state;
    end
    if (metaReset) begin
      _T_2906 <= 9'h0;
    end else if (reset) begin
      _T_2906 <= 9'h0;
    end else if (_T_2898) begin
      if (c_first) begin
        if (tl_out__c_bits_opcode[0]) begin
          _T_2906 <= _T_2903;
        end else begin
          _T_2906 <= 9'h0;
        end
      end else begin
        _T_2906 <= _T_2908;
      end
    end
    if (metaReset) begin
      s2_release_data_valid <= 1'h0;
    end else begin
      s2_release_data_valid <= s1_release_data_valid & ~releaseRejected;
    end
    if (metaReset) begin
      s1_req_cmd <= 5'h0;
    end else if (s0_clk_en) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if (metaReset) begin
      s2_req_cmd <= 5'h0;
    end else if (_T_2761) begin
      if (grantIsCached) begin
        if (_T_390) begin
          s2_req_cmd <= s1_req_cmd;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_cmd <= 5'h0;
        end else if (_T_390) begin
          s2_req_cmd <= s1_req_cmd;
        end
      end else if (_T_390) begin
        s2_req_cmd <= s1_req_cmd;
      end
    end else if (_T_390) begin
      s2_req_cmd <= s1_req_cmd;
    end
    if (metaReset) begin
      pstore1_held <= 1'h0;
    end else begin
      pstore1_held <= _T_1058 & ~pstore_drain;
    end
    if (metaReset) begin
      pstore1_addr <= 40'h0;
    end else if (_T_887) begin
      pstore1_addr <= s1_req_addr;
    end
    if (metaReset) begin
      s1_req_addr <= 40'h0;
    end else if (s0_clk_en) begin
      s1_req_addr <= s0_req_addr;
    end
    if (metaReset) begin
      pstore1_mask <= 8'h0;
    end else if (_T_887) begin
      if (_T_53) begin
        pstore1_mask <= 8'h0;
      end else begin
        pstore1_mask <= s1_mask_xwr;
      end
    end
    if (metaReset) begin
      s1_req_size <= 2'h0;
    end else if (s0_clk_en) begin
      s1_req_size <= io_cpu_req_bits_size;
    end
    if (metaReset) begin
      pstore2_valid <= 1'h0;
    end else begin
      pstore2_valid <= _T_1064 | advance_pstore1;
    end
    if (metaReset) begin
      pstore2_addr <= 40'h0;
    end else if (advance_pstore1) begin
      pstore2_addr <= pstore1_addr;
    end
    if (metaReset) begin
      mask <= 8'h0;
    end else if (advance_pstore1) begin
      mask <= pstore1_mask[7:0];
    end
    if (metaReset) begin
      s2_not_nacked_in_s1 <= 1'h0;
    end else begin
      s2_not_nacked_in_s1 <= ~s1_nack;
    end
    if (metaReset) begin
      s2_hit_state_state <= 2'h0;
    end else if (_T_390) begin
      s2_hit_state_state <= s1_meta_hit_state_state;
    end
    if (metaReset) begin
      s1_req_tag <= 7'h0;
    end else if (s0_clk_en) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if (metaReset) begin
      s1_req_signed <= 1'h0;
    end else if (s0_clk_en) begin
      s1_req_signed <= io_cpu_req_bits_signed;
    end
    if (metaReset) begin
      s1_tlb_req_vaddr <= 40'h0;
    end else if (s0_clk_en) begin
      s1_tlb_req_vaddr <= s0_req_addr;
    end
    if (metaReset) begin
      s1_tlb_req_passthrough <= 1'h0;
    end else if (s0_clk_en) begin
      s1_tlb_req_passthrough <= s0_req_phys;
    end
    if (metaReset) begin
      s1_tlb_req_size <= 2'h0;
    end else if (s0_clk_en) begin
      s1_tlb_req_size <= io_cpu_req_bits_size;
    end
    if (metaReset) begin
      s1_tlb_req_cmd <= 5'h0;
    end else if (s0_clk_en) begin
      s1_tlb_req_cmd <= io_cpu_req_bits_cmd;
    end
    if (metaReset) begin
      s1_flush_valid <= 1'h0;
    end else begin
      s1_flush_valid <= _T_3109 & ~release_ack_wait;
    end
    if (metaReset) begin
      cached_grant_wait <= 1'h0;
    end else if (reset) begin
      cached_grant_wait <= 1'h0;
    end else if (_T_2761) begin
      if (grantIsCached) begin
        if (d_last) begin
          cached_grant_wait <= 1'h0;
        end else if (_T_2700) begin
          if (!(s2_uncached)) begin
            cached_grant_wait <= 1'h1;
          end
        end
      end else if (_T_2700) begin
        if (!(s2_uncached)) begin
          cached_grant_wait <= 1'h1;
        end
      end
    end else if (_T_2700) begin
      if (!(s2_uncached)) begin
        cached_grant_wait <= 1'h1;
      end
    end
    if (metaReset) begin
      uncachedInFlight_0 <= 1'h0;
    end else if (reset) begin
      uncachedInFlight_0 <= 1'h0;
    end else if (_T_2761) begin
      if (grantIsCached) begin
        if (_T_2700) begin
          if (s2_uncached) begin
            uncachedInFlight_0 <= _GEN_143;
          end
        end
      end else if (grantIsUncached) begin
        if (_T_2766) begin
          uncachedInFlight_0 <= 1'h0;
        end else if (_T_2700) begin
          if (s2_uncached) begin
            uncachedInFlight_0 <= _GEN_143;
          end
        end
      end else if (_T_2700) begin
        if (s2_uncached) begin
          uncachedInFlight_0 <= _GEN_143;
        end
      end
    end else if (_T_2700) begin
      if (s2_uncached) begin
        uncachedInFlight_0 <= _GEN_143;
      end
    end
    if (metaReset) begin
      uncachedReqs_0_addr <= 40'h0;
    end else if (_T_2700) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_addr <= s2_req_addr;
        end
      end
    end
    if (metaReset) begin
      uncachedReqs_0_tag <= 7'h0;
    end else if (_T_2700) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_tag <= s2_req_tag;
        end
      end
    end
    if (metaReset) begin
      uncachedReqs_0_size <= 2'h0;
    end else if (_T_2700) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_size <= s2_req_size;
        end
      end
    end
    if (metaReset) begin
      uncachedReqs_0_signed <= 1'h0;
    end else if (_T_2700) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_signed <= s2_req_signed;
        end
      end
    end
    if (metaReset) begin
      s1_did_read <= 1'h0;
    end else if (s0_clk_en) begin
      s1_did_read <= _T_224;
    end
    if (metaReset) begin
      s2_hit_way <= 4'h0;
    end else if (s1_valid_not_nacked) begin
      s2_hit_way <= s1_meta_hit_way;
    end
    if (metaReset) begin
      _T_672 <= 2'h0;
    end else if (_T_390) begin
      _T_672 <= s1_victim_way;
    end
    if (metaReset) begin
      s2_probe_way <= 4'h0;
    end else if (s1_probe) begin
      s2_probe_way <= s1_meta_hit_way;
    end
    if (metaReset) begin
      s2_req_addr <= 40'h0;
    end else if (_T_2761) begin
      if (grantIsCached) begin
        if (_T_390) begin
          s2_req_addr <= {{8'd0}, s1_paddr};
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_addr <= {{8'd0}, _T_2773};
        end else if (_T_390) begin
          s2_req_addr <= {{8'd0}, s1_paddr};
        end
      end else if (_T_390) begin
        s2_req_addr <= {{8'd0}, s1_paddr};
      end
    end else if (_T_390) begin
      s2_req_addr <= {{8'd0}, s1_paddr};
    end
    if (metaReset) begin
      s2_req_tag <= 7'h0;
    end else if (_T_2761) begin
      if (grantIsCached) begin
        if (_T_390) begin
          s2_req_tag <= s1_req_tag;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_tag <= uncachedReqs_0_tag;
        end else if (_T_390) begin
          s2_req_tag <= s1_req_tag;
        end
      end else if (_T_390) begin
        s2_req_tag <= s1_req_tag;
      end
    end else if (_T_390) begin
      s2_req_tag <= s1_req_tag;
    end
    if (metaReset) begin
      s2_req_size <= 2'h0;
    end else if (_T_2761) begin
      if (grantIsCached) begin
        if (_T_390) begin
          s2_req_size <= s1_req_size;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_size <= uncachedReqs_0_size;
        end else if (_T_390) begin
          s2_req_size <= s1_req_size;
        end
      end else if (_T_390) begin
        s2_req_size <= s1_req_size;
      end
    end else if (_T_390) begin
      s2_req_size <= s1_req_size;
    end
    if (metaReset) begin
      s2_req_signed <= 1'h0;
    end else if (_T_2761) begin
      if (grantIsCached) begin
        if (_T_390) begin
          s2_req_signed <= s1_req_signed;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_signed <= uncachedReqs_0_signed;
        end else if (_T_390) begin
          s2_req_signed <= s1_req_signed;
        end
      end else if (_T_390) begin
        s2_req_signed <= s1_req_signed;
      end
    end else if (_T_390) begin
      s2_req_signed <= s1_req_signed;
    end
    if (metaReset) begin
      s2_tlb_xcpt_pf_ld <= 1'h0;
    end else if (_T_390) begin
      s2_tlb_xcpt_pf_ld <= tlb_io_resp_pf_ld;
    end
    if (metaReset) begin
      s2_tlb_xcpt_pf_st <= 1'h0;
    end else if (_T_390) begin
      s2_tlb_xcpt_pf_st <= tlb_io_resp_pf_st;
    end
    if (metaReset) begin
      s2_tlb_xcpt_ae_ld <= 1'h0;
    end else if (_T_390) begin
      s2_tlb_xcpt_ae_ld <= tlb_io_resp_ae_ld;
    end
    if (metaReset) begin
      s2_tlb_xcpt_ae_st <= 1'h0;
    end else if (_T_390) begin
      s2_tlb_xcpt_ae_st <= tlb_io_resp_ae_st;
    end
    if (metaReset) begin
      s2_tlb_xcpt_ma_ld <= 1'h0;
    end else if (_T_390) begin
      s2_tlb_xcpt_ma_ld <= tlb_io_resp_ma_ld;
    end
    if (metaReset) begin
      s2_tlb_xcpt_ma_st <= 1'h0;
    end else if (_T_390) begin
      s2_tlb_xcpt_ma_st <= tlb_io_resp_ma_st;
    end
    if (metaReset) begin
      s2_pma_cacheable <= 1'h0;
    end else if (_T_390) begin
      s2_pma_cacheable <= _T_391_cacheable;
    end
    if (metaReset) begin
      _T_393 <= 40'h0;
    end else if (_T_390) begin
      _T_393 <= s1_req_addr;
    end
    if (metaReset) begin
      s2_flush_valid_pre_tag_ecc <= 1'h0;
    end else begin
      s2_flush_valid_pre_tag_ecc <= s1_flush_valid;
    end
    if (metaReset) begin
      _T_465 <= 22'h0;
    end else if (s1_meta_clk_en) begin
      _T_465 <= tag_array_3_s1_meta_data;
    end
    if (metaReset) begin
      blockUncachedGrant <= 1'h0;
    end else if (_T_2878) begin
      if (auto_out_d_valid) begin
        blockUncachedGrant <= ~dataArb_io_in_1_ready;
      end else begin
        blockUncachedGrant <= dataArb_io_out_valid;
      end
    end else begin
      blockUncachedGrant <= dataArb_io_out_valid;
    end
    if (metaReset) begin
      _T_2713 <= 9'h0;
    end else if (reset) begin
      _T_2713 <= 9'h0;
    end else if (_T_2761) begin
      if (d_first) begin
        if (auto_out_d_bits_opcode[0]) begin
          _T_2713 <= _T_2710;
        end else begin
          _T_2713 <= 9'h0;
        end
      end else begin
        _T_2713 <= _T_2715;
      end
    end
    if (metaReset) begin
      s2_data <= 64'h0;
    end else if (en) begin
      s2_data <= _T_490;
    end
    if (metaReset) begin
      _T_677 <= 20'h0;
    end else if (_T_390) begin
      if (_T_320) begin
        _T_677 <= s1_meta_uncorrected_3_tag;
      end else if (_T_318) begin
        _T_677 <= s1_meta_uncorrected_2_tag;
      end else if (_T_316) begin
        _T_677 <= s1_meta_uncorrected_1_tag;
      end else begin
        _T_677 <= s1_meta_uncorrected_0_tag;
      end
    end
    if (metaReset) begin
      _T_679_state <= 2'h0;
    end else if (_T_390) begin
      if (_T_320) begin
        _T_679_state <= s1_meta_uncorrected_3_coh_state;
      end else if (_T_318) begin
        _T_679_state <= s1_meta_uncorrected_2_coh_state;
      end else if (_T_316) begin
        _T_679_state <= s1_meta_uncorrected_1_coh_state;
      end else begin
        _T_679_state <= s1_meta_uncorrected_0_coh_state;
      end
    end
    if (metaReset) begin
      lrscAddr <= 34'h0;
    end else if (_T_871) begin
      lrscAddr <= s2_req_addr[39:6];
    end
    if (metaReset) begin
      pstore1_cmd <= 5'h0;
    end else if (_T_887) begin
      pstore1_cmd <= s1_req_cmd;
    end
    if (metaReset) begin
      pstore1_data <= 64'h0;
    end else if (_T_887) begin
      pstore1_data <= io_cpu_s1_data_data;
    end
    if (metaReset) begin
      pstore1_way <= 4'h0;
    end else if (_T_887) begin
      pstore1_way <= s1_meta_hit_way;
    end
    if (metaReset) begin
      pstore1_rmw <= 1'h0;
    end else if (_T_887) begin
      pstore1_rmw <= _T_942;
    end
    if (metaReset) begin
      _T_1016 <= 1'h0;
    end else begin
      _T_1016 <= io_cpu_s2_nack;
    end
    if (metaReset) begin
      pstore2_way <= 4'h0;
    end else if (advance_pstore1) begin
      pstore2_way <= pstore1_way;
    end
    if (metaReset) begin
      _T_1072 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1072 <= pstore1_storegen_data[7:0];
    end
    if (metaReset) begin
      _T_1077 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1077 <= pstore1_storegen_data[15:8];
    end
    if (metaReset) begin
      _T_1082 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1082 <= pstore1_storegen_data[23:16];
    end
    if (metaReset) begin
      _T_1087 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1087 <= pstore1_storegen_data[31:24];
    end
    if (metaReset) begin
      _T_1092 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1092 <= pstore1_storegen_data[39:32];
    end
    if (metaReset) begin
      _T_1097 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1097 <= pstore1_storegen_data[47:40];
    end
    if (metaReset) begin
      _T_1102 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1102 <= pstore1_storegen_data[55:48];
    end
    if (metaReset) begin
      _T_1107 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1107 <= pstore1_storegen_data[63:56];
    end
    if (metaReset) begin
      s1_release_data_valid <= 1'h0;
    end else begin
      s1_release_data_valid <= dataArb_io_in_2_ready & dataArb_io_in_2_valid;
    end
    if (metaReset) begin
      _T_3014 <= 1'h0;
    end else begin
      _T_3014 <= _T_3012 & ~s1_nack;
    end
    if (metaReset) begin
      doUncachedResp <= 1'h0;
    end else begin
      doUncachedResp <= io_cpu_replay_next;
    end
    if (metaReset) begin
      resetting <= 1'h0;
    end else if (reset) begin
      resetting <= 1'h0;
    end else if (resetting) begin
      if (flushDone) begin
        resetting <= 1'h0;
      end else begin
        resetting <= _GEN_341;
      end
    end else begin
      resetting <= _GEN_341;
    end
    if (metaReset) begin
      _T_3097 <= 1'h0;
    end else begin
      _T_3097 <= reset;
    end
    if (metaReset) begin
      flushCounter <= 8'h0;
    end else if (reset) begin
      flushCounter <= 8'hc0;
    end else begin
      flushCounter <= _GEN_343[7:0];
    end
    if (metaReset) begin
      _T_3178 <= 9'h0;
    end else if (reset) begin
      _T_3178 <= 9'h0;
    end else if (_T_2898) begin
      if (_T_3181) begin
        if (tl_out__c_bits_opcode[0]) begin
          _T_3178 <= _T_2903;
        end else begin
          _T_3178 <= 9'h0;
        end
      end else begin
        _T_3178 <= _T_3180;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_165) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:1081 assert(!needsRead(req) || res)\n"); // @[DCache.scala 1081:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_165) begin
          $fatal; // @[DCache.scala 1081:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_370) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:281 assert(!(s1_valid_masked && s1_req.cmd === M_PWR) || (s1_mask_xwr | ~io.cpu.s1_data.mask).andR)\n"); // @[DCache.scala 281:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_370) begin
          $fatal; // @[DCache.scala 281:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_165) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:1081 assert(!needsRead(req) || res)\n"); // @[DCache.scala 1081:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_165) begin
          $fatal; // @[DCache.scala 1081:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1034) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:461 assert(pstore1_rmw || pstore1_valid_not_rmw(io.cpu.s2_kill) === pstore1_valid)\n"); // @[DCache.scala 461:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1034) begin
          $fatal; // @[DCache.scala 461:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_356 & ~_T_2763) begin
          $fwrite(32'h80000002,"Assertion failed: A GrantData was unexpected by the dcache.\n    at DCache.scala:620 assert(cached_grant_wait, \"A GrantData was unexpected by the dcache.\")\n"); // @[DCache.scala 620:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_356 & ~_T_2763) begin
          $fatal; // @[DCache.scala 620:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & ~_T_2768) begin
          $fwrite(32'h80000002,"Assertion failed: An AccessAck was unexpected by the dcache.\n    at DCache.scala:630 assert(f, \"An AccessAck was unexpected by the dcache.\") // TODO must handle Ack coming back on same cycle!\n"); // @[DCache.scala 630:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & ~_T_2768) begin
          $fatal; // @[DCache.scala 630:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_370 & ~_T_2775) begin
          $fwrite(32'h80000002,"Assertion failed: A ReleaseAck was unexpected by the dcache.\n    at DCache.scala:651 assert(release_ack_wait, \"A ReleaseAck was unexpected by the dcache.\") // TODO should handle Ack coming back on same cycle!\n"); // @[DCache.scala 651:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_370 & ~_T_2775) begin
          $fatal; // @[DCache.scala 651:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_2787) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:659 assert(tl_out.e.fire() === (tl_out.d.fire() && d_first && grantIsCached))\n"); // @[DCache.scala 659:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2787) begin
          $fatal; // @[DCache.scala 659:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s2_want_victimize & ~_T_2931) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:739 assert(s2_valid_flush_line || s2_flush_valid || io.cpu.s2_nack)\n"); // @[DCache.scala 739:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (s2_want_victimize & ~_T_2931) begin
          $fatal; // @[DCache.scala 739:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doUncachedResp & ~_T_3027) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:851 assert(!s2_valid_hit)\n"); // @[DCache.scala 851:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doUncachedResp & ~_T_3027) begin
          $fatal; // @[DCache.scala 851:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    DCache_state <= DCache_xor0;
    if (!(DCache_cov_read_data)) begin
      DCache_covSum <= DCache_covSum + 1'h1;
    end
  end
  always @(posedge gated_clock) begin
    if(DCache_cov_write_en & DCache_cov_write_mask) begin
      DCache_cov[DCache_cov_write_addr] <= DCache_cov_write_data; // @[Coverage map for DCache]
    end
  end
endmodule
module Frontend(
  input         gated_clock,
  input         reset,
  input         auto_icache_master_out_a_ready,
  output        auto_icache_master_out_a_valid,
  output [31:0] auto_icache_master_out_a_bits_address,
  input         auto_icache_master_out_d_valid,
  input  [2:0]  auto_icache_master_out_d_bits_opcode,
  input  [3:0]  auto_icache_master_out_d_bits_size,
  input  [63:0] auto_icache_master_out_d_bits_data,
  input         auto_icache_master_out_d_bits_corrupt,
  input  [31:0] auto_reset_vector_sink_in,
  input         io_cpu_might_request,
  input         io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_pc,
  input         io_cpu_req_bits_speculative,
  input         io_cpu_sfence_valid,
  input         io_cpu_sfence_bits_rs1,
  input         io_cpu_sfence_bits_rs2,
  input  [38:0] io_cpu_sfence_bits_addr,
  input         io_cpu_resp_ready,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_btb_taken,
  output        io_cpu_resp_bits_btb_bridx,
  output [4:0]  io_cpu_resp_bits_btb_entry,
  output [7:0]  io_cpu_resp_bits_btb_bht_history,
  output [39:0] io_cpu_resp_bits_pc,
  output [31:0] io_cpu_resp_bits_data,
  output        io_cpu_resp_bits_xcpt_pf_inst,
  output        io_cpu_resp_bits_xcpt_ae_inst,
  output        io_cpu_resp_bits_replay,
  input         io_cpu_btb_update_valid,
  input  [4:0]  io_cpu_btb_update_bits_prediction_entry,
  input  [38:0] io_cpu_btb_update_bits_pc,
  input         io_cpu_btb_update_bits_isValid,
  input  [38:0] io_cpu_btb_update_bits_br_pc,
  input  [1:0]  io_cpu_btb_update_bits_cfiType,
  input         io_cpu_bht_update_valid,
  input  [7:0]  io_cpu_bht_update_bits_prediction_history,
  input  [38:0] io_cpu_bht_update_bits_pc,
  input         io_cpu_bht_update_bits_branch,
  input         io_cpu_bht_update_bits_taken,
  input         io_cpu_bht_update_bits_mispredict,
  input         io_cpu_flush_icache,
  output [39:0] io_cpu_npc,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output        io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input         io_ptw_status_debug,
  input  [1:0]  io_ptw_status_prv,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input  [63:0] io_ptw_customCSRs_csrs_0_value,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         icache_halt,
  input         fq_halt,
  input         tlb_halt,
  input         btb_halt,
output [5:0]	 Checking_Frontend_regstate,	//Jaewon_regstate
  output [29:0]	 Checking_Frontend_covSum,	//Jaewon_regstate
    output [63:0]	 Checking_Frontend_covmap	//Jaewon_regstate
    );
      assign Checking_Frontend_regstate = Frontend_state;		//Jaewon_regstate
        assign Checking_Frontend_covSum = Frontend_covSum;		//Jaewon_regstate
	  assign Checking_Frontend_covmap = {Frontend_cov[0],Frontend_cov[1],Frontend_cov[2],Frontend_cov[3],Frontend_cov[4],Frontend_cov[5],Frontend_cov[6],Frontend_cov[7],Frontend_cov[8],Frontend_cov[9],  Frontend_cov[10],Frontend_cov[11],Frontend_cov[12],Frontend_cov[13],Frontend_cov[14],  Frontend_cov[15],Frontend_cov[16],Frontend_cov[17],Frontend_cov[18],Frontend_cov[19],Frontend_cov[20],Frontend_cov[21],Frontend_cov[22],Frontend_cov[23],Frontend_cov[24],Frontend_cov[25],Frontend_cov[26],Frontend_cov[27],Frontend_cov[28],Frontend_cov[29],Frontend_cov[30],Frontend_cov[31],Frontend_cov[32],Frontend_cov[33],Frontend_cov[34],   Frontend_cov[35],Frontend_cov[36],Frontend_cov[37],Frontend_cov[38],Frontend_cov[39],Frontend_cov[40],	Frontend_cov[41],Frontend_cov[42],Frontend_cov[43],Frontend_cov[44],   Frontend_cov[45],Frontend_cov[46],Frontend_cov[47],Frontend_cov[48],Frontend_cov[49],Frontend_cov[50],	Frontend_cov[51],Frontend_cov[52],Frontend_cov[53],Frontend_cov[54],  Frontend_cov[55],Frontend_cov[56],Frontend_cov[57],Frontend_cov[58],Frontend_cov[59],Frontend_cov[60],Frontend_cov[61],Frontend_cov[62],Frontend_cov[63]};		//Jaewon_regstate
  wire  icache_clock; // @[Frontend.scala 64:26]
  wire  icache_reset; // @[Frontend.scala 64:26]
  wire  icache_auto_master_out_a_ready; // @[Frontend.scala 64:26]
  wire  icache_auto_master_out_a_valid; // @[Frontend.scala 64:26]
  wire [31:0] icache_auto_master_out_a_bits_address; // @[Frontend.scala 64:26]
  wire  icache_auto_master_out_d_valid; // @[Frontend.scala 64:26]
  wire [2:0] icache_auto_master_out_d_bits_opcode; // @[Frontend.scala 64:26]
  wire [3:0] icache_auto_master_out_d_bits_size; // @[Frontend.scala 64:26]
  wire [63:0] icache_auto_master_out_d_bits_data; // @[Frontend.scala 64:26]
  wire  icache_auto_master_out_d_bits_corrupt; // @[Frontend.scala 64:26]
  wire  icache_io_req_ready; // @[Frontend.scala 64:26]
  wire  icache_io_req_valid; // @[Frontend.scala 64:26]
  wire [38:0] icache_io_req_bits_addr; // @[Frontend.scala 64:26]
  wire [31:0] icache_io_s1_paddr; // @[Frontend.scala 64:26]
  wire  icache_io_s1_kill; // @[Frontend.scala 64:26]
  wire  icache_io_s2_kill; // @[Frontend.scala 64:26]
  wire  icache_io_resp_valid; // @[Frontend.scala 64:26]
  wire [31:0] icache_io_resp_bits_data; // @[Frontend.scala 64:26]
  wire  icache_io_resp_bits_replay; // @[Frontend.scala 64:26]
  wire  icache_io_resp_bits_ae; // @[Frontend.scala 64:26]
  wire  icache_io_invalidate; // @[Frontend.scala 64:26]
  wire [29:0] icache_io_covSum; // @[Frontend.scala 64:26]
  wire  icache_metaAssert; // @[Frontend.scala 64:26]
  wire  icache_metaReset; // @[Frontend.scala 64:26]
  wire  icache_MaxPeriodFibonacciLFSR_halt; // @[Frontend.scala 64:26]
  wire  fq_clock; // @[Frontend.scala 86:57]
  wire  fq_reset; // @[Frontend.scala 86:57]
  wire  fq_io_enq_ready; // @[Frontend.scala 86:57]
  wire  fq_io_enq_valid; // @[Frontend.scala 86:57]
  wire  fq_io_enq_bits_btb_taken; // @[Frontend.scala 86:57]
  wire  fq_io_enq_bits_btb_bridx; // @[Frontend.scala 86:57]
  wire [4:0] fq_io_enq_bits_btb_entry; // @[Frontend.scala 86:57]
  wire [7:0] fq_io_enq_bits_btb_bht_history; // @[Frontend.scala 86:57]
  wire [39:0] fq_io_enq_bits_pc; // @[Frontend.scala 86:57]
  wire [31:0] fq_io_enq_bits_data; // @[Frontend.scala 86:57]
  wire [1:0] fq_io_enq_bits_mask; // @[Frontend.scala 86:57]
  wire  fq_io_enq_bits_xcpt_pf_inst; // @[Frontend.scala 86:57]
  wire  fq_io_enq_bits_xcpt_ae_inst; // @[Frontend.scala 86:57]
  wire  fq_io_enq_bits_replay; // @[Frontend.scala 86:57]
  wire  fq_io_deq_ready; // @[Frontend.scala 86:57]
  wire  fq_io_deq_valid; // @[Frontend.scala 86:57]
  wire  fq_io_deq_bits_btb_taken; // @[Frontend.scala 86:57]
  wire  fq_io_deq_bits_btb_bridx; // @[Frontend.scala 86:57]
  wire [4:0] fq_io_deq_bits_btb_entry; // @[Frontend.scala 86:57]
  wire [7:0] fq_io_deq_bits_btb_bht_history; // @[Frontend.scala 86:57]
  wire [39:0] fq_io_deq_bits_pc; // @[Frontend.scala 86:57]
  wire [31:0] fq_io_deq_bits_data; // @[Frontend.scala 86:57]
  wire  fq_io_deq_bits_xcpt_pf_inst; // @[Frontend.scala 86:57]
  wire  fq_io_deq_bits_xcpt_ae_inst; // @[Frontend.scala 86:57]
  wire  fq_io_deq_bits_replay; // @[Frontend.scala 86:57]
  wire [4:0] fq_io_mask; // @[Frontend.scala 86:57]
  wire [29:0] fq_io_covSum; // @[Frontend.scala 86:57]
  wire  fq_metaAssert; // @[Frontend.scala 86:57]
  wire  fq_metaReset; // @[Frontend.scala 86:57]
  wire  tlb_clock; // @[Frontend.scala 100:19]
  wire  tlb_reset; // @[Frontend.scala 100:19]
  wire  tlb_io_req_ready; // @[Frontend.scala 100:19]
  wire  tlb_io_req_valid; // @[Frontend.scala 100:19]
  wire [39:0] tlb_io_req_bits_vaddr; // @[Frontend.scala 100:19]
  wire  tlb_io_resp_miss; // @[Frontend.scala 100:19]
  wire [31:0] tlb_io_resp_paddr; // @[Frontend.scala 100:19]
  wire  tlb_io_resp_pf_inst; // @[Frontend.scala 100:19]
  wire  tlb_io_resp_ae_inst; // @[Frontend.scala 100:19]
  wire  tlb_io_resp_cacheable; // @[Frontend.scala 100:19]
  wire  tlb_io_sfence_valid; // @[Frontend.scala 100:19]
  wire  tlb_io_sfence_bits_rs1; // @[Frontend.scala 100:19]
  wire  tlb_io_sfence_bits_rs2; // @[Frontend.scala 100:19]
  wire [38:0] tlb_io_sfence_bits_addr; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_req_ready; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_req_valid; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_req_bits_valid; // @[Frontend.scala 100:19]
  wire [26:0] tlb_io_ptw_req_bits_bits_addr; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_resp_valid; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_resp_bits_ae; // @[Frontend.scala 100:19]
  wire [53:0] tlb_io_ptw_resp_bits_pte_ppn; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_resp_bits_pte_d; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_resp_bits_pte_a; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_resp_bits_pte_g; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_resp_bits_pte_u; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_resp_bits_pte_x; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_resp_bits_pte_w; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_resp_bits_pte_r; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_resp_bits_pte_v; // @[Frontend.scala 100:19]
  wire [1:0] tlb_io_ptw_resp_bits_level; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_resp_bits_homogeneous; // @[Frontend.scala 100:19]
  wire [3:0] tlb_io_ptw_ptbr_mode; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_status_debug; // @[Frontend.scala 100:19]
  wire [1:0] tlb_io_ptw_status_prv; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_0_cfg_l; // @[Frontend.scala 100:19]
  wire [1:0] tlb_io_ptw_pmp_0_cfg_a; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_0_cfg_x; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_0_cfg_w; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_0_cfg_r; // @[Frontend.scala 100:19]
  wire [29:0] tlb_io_ptw_pmp_0_addr; // @[Frontend.scala 100:19]
  wire [31:0] tlb_io_ptw_pmp_0_mask; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_1_cfg_l; // @[Frontend.scala 100:19]
  wire [1:0] tlb_io_ptw_pmp_1_cfg_a; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_1_cfg_x; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_1_cfg_w; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_1_cfg_r; // @[Frontend.scala 100:19]
  wire [29:0] tlb_io_ptw_pmp_1_addr; // @[Frontend.scala 100:19]
  wire [31:0] tlb_io_ptw_pmp_1_mask; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_2_cfg_l; // @[Frontend.scala 100:19]
  wire [1:0] tlb_io_ptw_pmp_2_cfg_a; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_2_cfg_x; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_2_cfg_w; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_2_cfg_r; // @[Frontend.scala 100:19]
  wire [29:0] tlb_io_ptw_pmp_2_addr; // @[Frontend.scala 100:19]
  wire [31:0] tlb_io_ptw_pmp_2_mask; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_3_cfg_l; // @[Frontend.scala 100:19]
  wire [1:0] tlb_io_ptw_pmp_3_cfg_a; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_3_cfg_x; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_3_cfg_w; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_3_cfg_r; // @[Frontend.scala 100:19]
  wire [29:0] tlb_io_ptw_pmp_3_addr; // @[Frontend.scala 100:19]
  wire [31:0] tlb_io_ptw_pmp_3_mask; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_4_cfg_l; // @[Frontend.scala 100:19]
  wire [1:0] tlb_io_ptw_pmp_4_cfg_a; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_4_cfg_x; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_4_cfg_w; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_4_cfg_r; // @[Frontend.scala 100:19]
  wire [29:0] tlb_io_ptw_pmp_4_addr; // @[Frontend.scala 100:19]
  wire [31:0] tlb_io_ptw_pmp_4_mask; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_5_cfg_l; // @[Frontend.scala 100:19]
  wire [1:0] tlb_io_ptw_pmp_5_cfg_a; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_5_cfg_x; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_5_cfg_w; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_5_cfg_r; // @[Frontend.scala 100:19]
  wire [29:0] tlb_io_ptw_pmp_5_addr; // @[Frontend.scala 100:19]
  wire [31:0] tlb_io_ptw_pmp_5_mask; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_6_cfg_l; // @[Frontend.scala 100:19]
  wire [1:0] tlb_io_ptw_pmp_6_cfg_a; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_6_cfg_x; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_6_cfg_w; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_6_cfg_r; // @[Frontend.scala 100:19]
  wire [29:0] tlb_io_ptw_pmp_6_addr; // @[Frontend.scala 100:19]
  wire [31:0] tlb_io_ptw_pmp_6_mask; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_7_cfg_l; // @[Frontend.scala 100:19]
  wire [1:0] tlb_io_ptw_pmp_7_cfg_a; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_7_cfg_x; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_7_cfg_w; // @[Frontend.scala 100:19]
  wire  tlb_io_ptw_pmp_7_cfg_r; // @[Frontend.scala 100:19]
  wire [29:0] tlb_io_ptw_pmp_7_addr; // @[Frontend.scala 100:19]
  wire [31:0] tlb_io_ptw_pmp_7_mask; // @[Frontend.scala 100:19]
  wire  tlb_io_kill; // @[Frontend.scala 100:19]
  wire [29:0] tlb_io_covSum; // @[Frontend.scala 100:19]
  wire  tlb_metaAssert; // @[Frontend.scala 100:19]
  wire  tlb_metaReset; // @[Frontend.scala 100:19]
  wire  btb_clock; // @[Frontend.scala 181:21]
  wire  btb_reset; // @[Frontend.scala 181:21]
  wire [38:0] btb_io_req_bits_addr; // @[Frontend.scala 181:21]
  wire  btb_io_resp_valid; // @[Frontend.scala 181:21]
  wire  btb_io_resp_bits_taken; // @[Frontend.scala 181:21]
  wire  btb_io_resp_bits_bridx; // @[Frontend.scala 181:21]
  wire [38:0] btb_io_resp_bits_target; // @[Frontend.scala 181:21]
  wire [4:0] btb_io_resp_bits_entry; // @[Frontend.scala 181:21]
  wire [7:0] btb_io_resp_bits_bht_history; // @[Frontend.scala 181:21]
  wire  btb_io_resp_bits_bht_value; // @[Frontend.scala 181:21]
  wire  btb_io_btb_update_valid; // @[Frontend.scala 181:21]
  wire [4:0] btb_io_btb_update_bits_prediction_entry; // @[Frontend.scala 181:21]
  wire [38:0] btb_io_btb_update_bits_pc; // @[Frontend.scala 181:21]
  wire  btb_io_btb_update_bits_isValid; // @[Frontend.scala 181:21]
  wire [38:0] btb_io_btb_update_bits_br_pc; // @[Frontend.scala 181:21]
  wire [1:0] btb_io_btb_update_bits_cfiType; // @[Frontend.scala 181:21]
  wire  btb_io_bht_update_valid; // @[Frontend.scala 181:21]
  wire [7:0] btb_io_bht_update_bits_prediction_history; // @[Frontend.scala 181:21]
  wire [38:0] btb_io_bht_update_bits_pc; // @[Frontend.scala 181:21]
  wire  btb_io_bht_update_bits_branch; // @[Frontend.scala 181:21]
  wire  btb_io_bht_update_bits_taken; // @[Frontend.scala 181:21]
  wire  btb_io_bht_update_bits_mispredict; // @[Frontend.scala 181:21]
  wire  btb_io_bht_advance_valid; // @[Frontend.scala 181:21]
  wire  btb_io_bht_advance_bits_bht_value; // @[Frontend.scala 181:21]
  wire  btb_io_ras_update_valid; // @[Frontend.scala 181:21]
  wire [1:0] btb_io_ras_update_bits_cfiType; // @[Frontend.scala 181:21]
  wire [38:0] btb_io_ras_update_bits_returnAddr; // @[Frontend.scala 181:21]
  wire  btb_io_ras_head_valid; // @[Frontend.scala 181:21]
  wire [38:0] btb_io_ras_head_bits; // @[Frontend.scala 181:21]
  wire  btb_io_flush; // @[Frontend.scala 181:21]
  wire [29:0] btb_io_covSum; // @[Frontend.scala 181:21]
  wire  btb_metaAssert; // @[Frontend.scala 181:21]
  wire  btb_metaReset; // @[Frontend.scala 181:21]
  wire  _T_2; // @[Frontend.scala 91:29]
  wire  _T_3; // @[Frontend.scala 91:52]
  wire  _T_4; // @[Frontend.scala 91:75]
  wire  _T_5; // @[Frontend.scala 91:102]
  wire  _T_7; // @[Frontend.scala 91:130]
  wire  _T_9; // @[Frontend.scala 91:9]
  reg  s1_valid; // @[Frontend.scala 102:21]
  reg [31:0] _RAND_0;
  reg  s2_valid; // @[Frontend.scala 103:25]
  reg [31:0] _RAND_1;
  wire  _T_17; // @[Frontend.scala 106:55]
  wire  _T_18; // @[Frontend.scala 106:41]
  wire  _T_19; // @[Frontend.scala 105:40]
  wire  _T_24; // @[Frontend.scala 107:55]
  wire  _T_25; // @[Frontend.scala 107:41]
  wire  s0_fq_has_space; // @[Frontend.scala 106:70]
  wire  s0_valid; // @[Frontend.scala 108:35]
  reg [39:0] s1_pc; // @[Frontend.scala 110:18]
  reg [63:0] _RAND_2;
  reg  s1_speculative; // @[Frontend.scala 111:27]
  reg [31:0] _RAND_3;
  wire [31:0] _T_27; // @[Frontend.scala 343:33]
  reg [39:0] s2_pc; // @[Frontend.scala 112:22]
  reg [63:0] _RAND_4;
  reg  s2_btb_resp_valid; // @[Frontend.scala 113:44]
  reg [31:0] _RAND_5;
  reg  s2_btb_resp_bits_taken; // @[Frontend.scala 114:29]
  reg [31:0] _RAND_6;
  reg  s2_btb_resp_bits_bridx; // @[Frontend.scala 114:29]
  reg [31:0] _RAND_7;
  reg [4:0] s2_btb_resp_bits_entry; // @[Frontend.scala 114:29]
  reg [31:0] _RAND_8;
  reg [7:0] s2_btb_resp_bits_bht_history; // @[Frontend.scala 114:29]
  reg [31:0] _RAND_9;
  reg  s2_btb_resp_bits_bht_value; // @[Frontend.scala 114:29]
  reg [31:0] _RAND_10;
  wire  s2_btb_taken; // @[Frontend.scala 115:40]
  reg  s2_tlb_resp_miss; // @[Frontend.scala 116:24]
  reg [31:0] _RAND_11;
  reg  s2_tlb_resp_pf_inst; // @[Frontend.scala 116:24]
  reg [31:0] _RAND_12;
  reg  s2_tlb_resp_ae_inst; // @[Frontend.scala 116:24]
  reg [31:0] _RAND_13;
  reg  s2_tlb_resp_cacheable; // @[Frontend.scala 116:24]
  reg [31:0] _RAND_14;
  wire  s2_xcpt; // @[Frontend.scala 117:37]
  reg  s2_speculative; // @[Frontend.scala 118:27]
  reg [31:0] _RAND_15;
  reg  s2_partial_insn_valid; // @[Frontend.scala 119:38]
  reg [31:0] _RAND_16;
  reg [15:0] s2_partial_insn; // @[Frontend.scala 120:28]
  reg [31:0] _RAND_17;
  reg  wrong_path; // @[Frontend.scala 121:23]
  reg [31:0] _RAND_18;
  wire [39:0] _T_30; // @[Frontend.scala 123:29]
  wire [39:0] s1_base_pc; // @[Frontend.scala 123:20]
  wire [39:0] ntpc; // @[Frontend.scala 124:25]
  wire  _T_32; // @[Decoupled.scala 40:37]
  wire  _T_34; // @[Frontend.scala 129:26]
  reg  _T_37; // @[Frontend.scala 129:58]
  reg [31:0] _RAND_19;
  wire  s2_replay; // @[Frontend.scala 129:48]
  wire  _T_36; // @[Frontend.scala 129:69]
  wire  _T_105; // @[Frontend.scala 210:45]
  wire  taken_prevRVI; // @[Frontend.scala 211:31]
  wire [15:0] taken_bits; // @[Frontend.scala 213:37]
  wire [31:0] taken_rviBits; // @[Cat.scala 29:58]
  wire  taken_rviJump; // @[Frontend.scala 217:34]
  wire  taken_rviJALR; // @[Frontend.scala 218:34]
  wire  _T_299; // @[Frontend.scala 232:29]
  wire  taken_rviBranch; // @[Frontend.scala 216:36]
  wire  _T_300; // @[Frontend.scala 232:53]
  wire  _T_301; // @[Frontend.scala 232:40]
  wire  _T_302; // @[Frontend.scala 232:17]
  wire  taken_valid; // @[Frontend.scala 212:44]
  wire [15:0] _T_127; // @[Frontend.scala 223:26]
  wire  taken_rvcJump; // @[Frontend.scala 223:26]
  wire [15:0] _T_169; // @[Frontend.scala 227:26]
  wire  _T_170; // @[Frontend.scala 227:26]
  wire  _T_172; // @[Frontend.scala 227:62]
  wire  taken_rvcJALR; // @[Frontend.scala 227:49]
  wire  _T_303; // @[Frontend.scala 233:27]
  wire  _T_163; // @[Frontend.scala 225:24]
  wire  taken_rvcJR; // @[Frontend.scala 225:46]
  wire  _T_304; // @[Frontend.scala 233:38]
  wire  _T_122; // @[Frontend.scala 221:28]
  wire  _T_124; // @[Frontend.scala 221:60]
  wire  taken_rvcBranch; // @[Frontend.scala 221:52]
  wire  _T_305; // @[Frontend.scala 233:60]
  wire  _T_306; // @[Frontend.scala 233:47]
  wire  _T_307; // @[Frontend.scala 233:15]
  wire  taken_taken; // @[Frontend.scala 232:71]
  wire  taken_idx; // @[Frontend.scala 247:13]
  wire  _T_372; // @[Frontend.scala 210:45]
  wire  taken_prevRVI_1; // @[Frontend.scala 211:31]
  wire [15:0] taken_bits_1; // @[Frontend.scala 213:37]
  wire [31:0] taken_rviBits_1; // @[Cat.scala 29:58]
  wire  taken_rviJALR_1; // @[Frontend.scala 218:34]
  wire  _T_382; // @[Frontend.scala 219:31]
  wire [4:0] _T_384; // @[Frontend.scala 219:66]
  wire  _T_385; // @[Frontend.scala 219:66]
  wire  taken_rviReturn_1; // @[Frontend.scala 219:46]
  wire  _T_575; // @[Frontend.scala 234:61]
  wire  taken_valid_1; // @[Frontend.scala 212:44]
  wire [15:0] _T_429; // @[Frontend.scala 225:24]
  wire  _T_430; // @[Frontend.scala 225:24]
  wire  _T_432; // @[Frontend.scala 225:59]
  wire  taken_rvcJR_1; // @[Frontend.scala 225:46]
  wire [4:0] _T_434; // @[Frontend.scala 226:49]
  wire  _T_435; // @[Frontend.scala 226:49]
  wire  taken_rvcReturn_1; // @[Frontend.scala 226:29]
  wire  _T_576; // @[Frontend.scala 234:83]
  wire  _T_577; // @[Frontend.scala 234:74]
  wire  taken_predictReturn_1; // @[Frontend.scala 234:49]
  wire  _T_616; // @[Frontend.scala 260:26]
  wire  _T_115; // @[Frontend.scala 219:31]
  wire [4:0] _T_117; // @[Frontend.scala 219:66]
  wire  _T_118; // @[Frontend.scala 219:66]
  wire  taken_rviReturn; // @[Frontend.scala 219:46]
  wire  _T_308; // @[Frontend.scala 234:61]
  wire [4:0] _T_167; // @[Frontend.scala 226:49]
  wire  _T_168; // @[Frontend.scala 226:49]
  wire  taken_rvcReturn; // @[Frontend.scala 226:29]
  wire  _T_309; // @[Frontend.scala 234:83]
  wire  _T_310; // @[Frontend.scala 234:74]
  wire  taken_predictReturn; // @[Frontend.scala 234:49]
  wire  _T_349; // @[Frontend.scala 260:26]
  wire  _GEN_45; // @[Frontend.scala 256:30]
  wire  _GEN_78; // @[Frontend.scala 260:44]
  wire  _GEN_81; // @[Frontend.scala 256:30]
  wire  useRAS; // @[Frontend.scala 247:25]
  wire  taken_rviBranch_1; // @[Frontend.scala 216:36]
  wire  _T_580; // @[Frontend.scala 236:53]
  wire [15:0] _T_388; // @[Frontend.scala 221:28]
  wire  _T_389; // @[Frontend.scala 221:28]
  wire  _T_391; // @[Frontend.scala 221:60]
  wire  taken_rvcBranch_1; // @[Frontend.scala 221:52]
  wire  _T_581; // @[Frontend.scala 236:75]
  wire  _T_582; // @[Frontend.scala 236:66]
  wire  taken_predictBranch_1; // @[Frontend.scala 236:41]
  wire  taken_rviJump_1; // @[Frontend.scala 217:34]
  wire  _T_578; // @[Frontend.scala 235:33]
  wire  taken_rvcJump_1; // @[Frontend.scala 223:26]
  wire  _T_579; // @[Frontend.scala 235:53]
  wire  taken_predictJump_1; // @[Frontend.scala 235:44]
  wire  _T_617; // @[Frontend.scala 263:44]
  wire  _T_618; // @[Frontend.scala 263:26]
  wire [39:0] _T_91; // @[Frontend.scala 203:31]
  wire [39:0] s2_base_pc; // @[Frontend.scala 203:22]
  wire [39:0] taken_pc_1; // @[Frontend.scala 264:33]
  wire [39:0] _T_620; // @[Frontend.scala 267:36]
  wire [39:0] _T_622; // @[Frontend.scala 267:57]
  wire  _T_443; // @[RocketCore.scala 1036:53]
  wire  _T_498; // @[Cat.scala 29:58]
  wire [10:0] _T_497; // @[Cat.scala 29:58]
  wire [7:0] _T_495; // @[Cat.scala 29:58]
  wire  _T_494; // @[Cat.scala 29:58]
  wire [31:0] _T_502; // @[RocketCore.scala 1050:53]
  wire [7:0] _T_557; // @[Cat.scala 29:58]
  wire  _T_556; // @[Cat.scala 29:58]
  wire [31:0] _T_564; // @[RocketCore.scala 1050:53]
  wire [31:0] taken_rviImm_1; // @[Frontend.scala 229:23]
  wire [4:0] _T_399; // @[Bitwise.scala 72:12]
  wire [12:0] _T_409; // @[Frontend.scala 224:66]
  wire [9:0] _T_412; // @[Bitwise.scala 72:12]
  wire [20:0] _T_428; // @[Frontend.scala 224:106]
  wire [20:0] taken_rvcImm_1; // @[Frontend.scala 224:23]
  wire [31:0] _T_623; // @[Frontend.scala 267:69]
  wire [39:0] _GEN_127; // @[Frontend.scala 267:64]
  wire [39:0] _T_626; // @[Frontend.scala 268:34]
  wire  _T_313; // @[Frontend.scala 236:53]
  wire  _T_314; // @[Frontend.scala 236:75]
  wire  _T_315; // @[Frontend.scala 236:66]
  wire  taken_predictBranch; // @[Frontend.scala 236:41]
  wire  _T_311; // @[Frontend.scala 235:33]
  wire  _T_312; // @[Frontend.scala 235:53]
  wire  taken_predictJump; // @[Frontend.scala 235:44]
  wire  _T_350; // @[Frontend.scala 263:44]
  wire  _T_351; // @[Frontend.scala 263:26]
  wire [39:0] _T_352; // @[Frontend.scala 266:32]
  wire  _T_176; // @[RocketCore.scala 1036:53]
  wire  _T_231; // @[Cat.scala 29:58]
  wire [10:0] _T_230; // @[Cat.scala 29:58]
  wire [7:0] _T_228; // @[Cat.scala 29:58]
  wire  _T_227; // @[Cat.scala 29:58]
  wire [31:0] _T_235; // @[RocketCore.scala 1050:53]
  wire [7:0] _T_290; // @[Cat.scala 29:58]
  wire  _T_289; // @[Cat.scala 29:58]
  wire [31:0] _T_297; // @[RocketCore.scala 1050:53]
  wire [31:0] taken_rviImm; // @[Frontend.scala 229:23]
  wire [32:0] _T_353; // @[Frontend.scala 266:61]
  wire [4:0] _T_132; // @[Bitwise.scala 72:12]
  wire [12:0] _T_142; // @[Frontend.scala 224:66]
  wire [9:0] _T_145; // @[Bitwise.scala 72:12]
  wire [20:0] _T_161; // @[Frontend.scala 224:106]
  wire [20:0] taken_rvcImm; // @[Frontend.scala 224:23]
  wire [32:0] _T_354; // @[Frontend.scala 266:44]
  wire [39:0] _GEN_128; // @[Frontend.scala 266:39]
  wire [39:0] _T_357; // @[Frontend.scala 268:34]
  wire  predicted_taken; // @[Frontend.scala 194:29]
  wire [39:0] _T_89; // @[Cat.scala 29:58]
  wire [39:0] _GEN_28; // @[Frontend.scala 194:56]
  wire [39:0] _GEN_43; // @[Frontend.scala 263:61]
  wire [39:0] _GEN_46; // @[Frontend.scala 256:30]
  wire [39:0] _GEN_79; // @[Frontend.scala 263:61]
  wire [39:0] _GEN_82; // @[Frontend.scala 256:30]
  wire [39:0] _GEN_99; // @[Frontend.scala 247:25]
  wire [39:0] predicted_npc; // @[Frontend.scala 307:19]
  wire [39:0] npc; // @[Frontend.scala 130:16]
  wire  _T_40; // @[Frontend.scala 136:53]
  wire  _T_41; // @[Frontend.scala 136:41]
  wire  s0_speculative; // @[Frontend.scala 136:72]
  wire  _T_566; // @[Frontend.scala 232:29]
  wire  _T_567; // @[Frontend.scala 232:53]
  wire  _T_568; // @[Frontend.scala 232:40]
  wire  _T_569; // @[Frontend.scala 232:17]
  wire  _T_437; // @[Frontend.scala 227:26]
  wire  taken_rvcJALR_1; // @[Frontend.scala 227:49]
  wire  _T_570; // @[Frontend.scala 233:27]
  wire  _T_571; // @[Frontend.scala 233:38]
  wire  _T_572; // @[Frontend.scala 233:60]
  wire  _T_573; // @[Frontend.scala 233:47]
  wire  _T_574; // @[Frontend.scala 233:15]
  wire  taken_taken_1; // @[Frontend.scala 232:71]
  wire  taken; // @[Frontend.scala 288:19]
  wire  _GEN_116; // @[Frontend.scala 318:33]
  wire  _GEN_120; // @[Frontend.scala 314:20]
  wire  s2_redirect; // @[Frontend.scala 313:26]
  wire  _GEN_0; // @[Frontend.scala 142:21]
  wire  _T_49; // @[Frontend.scala 162:36]
  wire  s2_can_speculatively_refill; // @[Frontend.scala 163:59]
  wire  _T_54; // @[Frontend.scala 164:39]
  reg  _T_59; // @[Frontend.scala 167:29]
  reg [31:0] _RAND_20;
  wire  _T_60; // @[Frontend.scala 167:40]
  wire  _T_62; // @[Frontend.scala 167:98]
  wire  _T_63; // @[Frontend.scala 167:77]
  wire [39:0] _T_65; // @[Frontend.scala 169:28]
  wire [39:0] _T_67; // @[Frontend.scala 343:33]
  wire [2:0] _T_70; // @[Frontend.scala 172:52]
  wire  _T_72; // @[Frontend.scala 173:76]
  wire  _T_74; // @[Frontend.scala 173:101]
  wire  _T_75; // @[Frontend.scala 173:55]
  wire  _T_77; // @[Frontend.scala 177:27]
  wire  _T_79; // @[Frontend.scala 177:110]
  wire  _T_82; // @[Frontend.scala 177:9]
  wire  _T_84; // @[Frontend.scala 178:30]
  wire  fetch_bubble_likely; // @[Frontend.scala 295:33]
  wire  _T_96; // @[Frontend.scala 296:51]
  wire  _T_97; // @[Frontend.scala 296:66]
  wire  _T_635; // @[Frontend.scala 275:52]
  wire  _T_636; // @[Frontend.scala 275:91]
  wire  _T_637; // @[Frontend.scala 275:106]
  wire  _T_638; // @[Frontend.scala 275:34]
  wire  _T_366; // @[Frontend.scala 275:52]
  wire  _T_367; // @[Frontend.scala 275:91]
  wire  _T_368; // @[Frontend.scala 275:106]
  wire  _T_369; // @[Frontend.scala 275:34]
  wire  _GEN_92; // @[Frontend.scala 275:125]
  wire  updateBTB; // @[Frontend.scala 247:25]
  wire  _T_98; // @[Frontend.scala 296:89]
  wire [1:0] _T_99; // @[Frontend.scala 300:63]
  wire [39:0] _GEN_129; // @[Frontend.scala 300:50]
  wire [39:0] _T_100; // @[Frontend.scala 300:50]
  wire [39:0] _GEN_36; // @[Frontend.scala 294:37]
  wire [39:0] _GEN_37; // @[Frontend.scala 294:37]
  wire [1:0] after_idx; // @[Frontend.scala 247:25]
  wire [2:0] _T_101; // @[Frontend.scala 304:66]
  wire [39:0] _GEN_130; // @[Frontend.scala 304:53]
  wire [39:0] _T_103; // @[Frontend.scala 304:53]
  wire  _T_119; // @[Frontend.scala 220:30]
  wire  taken_rviCall; // @[Frontend.scala 220:42]
  wire  _T_316; // @[Frontend.scala 238:22]
  wire  _T_318; // @[Frontend.scala 238:43]
  wire  _T_319; // @[Frontend.scala 238:77]
  wire  _T_321; // @[Frontend.scala 238:86]
  wire  _GEN_39; // @[Frontend.scala 238:95]
  wire  _GEN_40; // @[Frontend.scala 238:95]
  wire  _T_326; // @[Frontend.scala 250:92]
  wire  _T_327; // @[Frontend.scala 250:80]
  wire  _T_328; // @[Frontend.scala 250:127]
  wire  _T_329; // @[Frontend.scala 250:115]
  wire  _T_330; // @[Frontend.scala 250:106]
  wire  _T_331; // @[Frontend.scala 250:68]
  wire  _T_332; // @[Frontend.scala 251:50]
  wire  _T_333; // @[Frontend.scala 252:50]
  wire  _T_334; // @[Frontend.scala 253:50]
  wire  _T_337; // @[Frontend.scala 253:46]
  wire [1:0] _T_338; // @[Frontend.scala 252:46]
  wire [1:0] _T_339; // @[Frontend.scala 251:46]
  wire  _T_342; // @[Frontend.scala 257:34]
  wire  _T_344; // @[Frontend.scala 257:43]
  wire  _T_346; // @[Frontend.scala 257:61]
  wire  _T_348; // @[Frontend.scala 257:77]
  wire  _GEN_41; // @[Frontend.scala 257:96]
  wire  _GEN_44; // @[Frontend.scala 256:30]
  wire  _GEN_47; // @[Frontend.scala 271:59]
  wire  taken_rvc_1; // @[Frontend.scala 210:45]
  wire  _T_386; // @[Frontend.scala 220:30]
  wire  taken_rviCall_1; // @[Frontend.scala 220:42]
  wire  _T_585; // @[Frontend.scala 238:43]
  wire  _T_586; // @[Frontend.scala 238:77]
  wire  _T_588; // @[Frontend.scala 238:86]
  wire  _GEN_76; // @[Frontend.scala 238:95]
  wire  _T_593; // @[Frontend.scala 250:92]
  wire  _T_594; // @[Frontend.scala 250:80]
  wire  _T_595; // @[Frontend.scala 250:127]
  wire  _T_596; // @[Frontend.scala 250:115]
  wire  _T_597; // @[Frontend.scala 250:106]
  wire  _T_598; // @[Frontend.scala 250:68]
  wire  _T_599; // @[Frontend.scala 251:50]
  wire  _T_600; // @[Frontend.scala 252:50]
  wire  _T_601; // @[Frontend.scala 253:50]
  wire  _T_604; // @[Frontend.scala 253:46]
  wire [1:0] _T_605; // @[Frontend.scala 252:46]
  wire [1:0] _T_606; // @[Frontend.scala 251:46]
  wire  _T_609; // @[Frontend.scala 257:34]
  wire  _T_611; // @[Frontend.scala 257:43]
  wire  _T_613; // @[Frontend.scala 257:61]
  wire  _T_615; // @[Frontend.scala 257:77]
  wire  _GEN_77; // @[Frontend.scala 257:96]
  wire  _GEN_83; // @[Frontend.scala 271:59]
  wire  _T_641; // @[Frontend.scala 283:23]
  wire  _T_643; // @[Frontend.scala 283:37]
  wire [15:0] _T_644; // @[Frontend.scala 285:37]
  wire  _T_646; // @[Frontend.scala 310:45]
  wire  _T_647; // @[Frontend.scala 310:28]
  wire  _GEN_117; // @[Frontend.scala 314:20]
  wire  _GEN_118; // @[Frontend.scala 314:20]
  wire [4:0] _GEN_119; // @[Frontend.scala 314:20]
  wire  _T_652; // @[Frontend.scala 322:35]
  wire  _T_654; // @[Frontend.scala 322:11]
  reg [5:0] Frontend_state; // @[Register tracking Frontend state]
  reg [31:0] _RAND_21;
  reg  Frontend_cov [0:63]; // @[Coverage map for Frontend]
  reg [31:0] _RAND_22;
  wire  Frontend_cov_read_data; // @[Coverage map for Frontend]
  wire [5:0] Frontend_cov_read_addr; // @[Coverage map for Frontend]
  wire  Frontend_cov_write_data; // @[Coverage map for Frontend]
  wire [5:0] Frontend_cov_write_addr; // @[Coverage map for Frontend]
  wire  Frontend_cov_write_mask; // @[Coverage map for Frontend]
  wire  Frontend_cov_write_en; // @[Coverage map for Frontend]
  reg [29:0] Frontend_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_23;
  wire  s2_partial_insn_valid_shl;
  wire [5:0] s2_partial_insn_valid_pad;
  wire [1:0] _T_37_shl;
  wire [5:0] _T_37_pad;
  wire [2:0] s2_btb_resp_valid_shl;
  wire [5:0] s2_btb_resp_valid_pad;
  wire [3:0] s2_btb_resp_bits_taken_shl;
  wire [5:0] s2_btb_resp_bits_taken_pad;
  wire [4:0] s2_btb_resp_bits_bht_value_shl;
  wire [5:0] s2_btb_resp_bits_bht_value_pad;
  wire [5:0] s2_valid_shl;
  wire [5:0] s2_valid_pad;
  wire [5:0] Frontend_xor4;
  wire [5:0] Frontend_xor1;
  wire [5:0] Frontend_xor6;
  wire [5:0] Frontend_xor2;
  wire [5:0] Frontend_xor0;
  wire [29:0] icache_sum;
  wire [29:0] fq_sum;
  wire [29:0] tlb_sum;
  wire [29:0] btb_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  icache_metaAssert_wire;
  wire  fq_metaAssert_wire;
  wire  tlb_metaAssert_wire;
  wire  btb_metaAssert_wire;
  wire  Frontend_or4;
  wire  Frontend_or1;
  wire  Frontend_or5;
  wire  Frontend_or6;
  wire  Frontend_or2;
  wire  Frontend_or0;
  ICache icache ( // @[Frontend.scala 64:26]
    .clock(icache_clock),
    .reset(icache_reset),
    .auto_master_out_a_ready(icache_auto_master_out_a_ready),
    .auto_master_out_a_valid(icache_auto_master_out_a_valid),
    .auto_master_out_a_bits_address(icache_auto_master_out_a_bits_address),
    .auto_master_out_d_valid(icache_auto_master_out_d_valid),
    .auto_master_out_d_bits_opcode(icache_auto_master_out_d_bits_opcode),
    .auto_master_out_d_bits_size(icache_auto_master_out_d_bits_size),
    .auto_master_out_d_bits_data(icache_auto_master_out_d_bits_data),
    .auto_master_out_d_bits_corrupt(icache_auto_master_out_d_bits_corrupt),
    .io_req_ready(icache_io_req_ready),
    .io_req_valid(icache_io_req_valid),
    .io_req_bits_addr(icache_io_req_bits_addr),
    .io_s1_paddr(icache_io_s1_paddr),
    .io_s1_kill(icache_io_s1_kill),
    .io_s2_kill(icache_io_s2_kill),
    .io_resp_valid(icache_io_resp_valid),
    .io_resp_bits_data(icache_io_resp_bits_data),
    .io_resp_bits_replay(icache_io_resp_bits_replay),
    .io_resp_bits_ae(icache_io_resp_bits_ae),
    .io_invalidate(icache_io_invalidate),
    .io_covSum(icache_io_covSum),
    .metaAssert(icache_metaAssert),
    .metaReset(icache_metaReset),
    .MaxPeriodFibonacciLFSR_halt(icache_MaxPeriodFibonacciLFSR_halt)
  );
  ShiftQueue fq ( // @[Frontend.scala 86:57]
    .clock(fq_clock),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_btb_taken(fq_io_enq_bits_btb_taken),
    .io_enq_bits_btb_bridx(fq_io_enq_bits_btb_bridx),
    .io_enq_bits_btb_entry(fq_io_enq_bits_btb_entry),
    .io_enq_bits_btb_bht_history(fq_io_enq_bits_btb_bht_history),
    .io_enq_bits_pc(fq_io_enq_bits_pc),
    .io_enq_bits_data(fq_io_enq_bits_data),
    .io_enq_bits_mask(fq_io_enq_bits_mask),
    .io_enq_bits_xcpt_pf_inst(fq_io_enq_bits_xcpt_pf_inst),
    .io_enq_bits_xcpt_ae_inst(fq_io_enq_bits_xcpt_ae_inst),
    .io_enq_bits_replay(fq_io_enq_bits_replay),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_btb_taken(fq_io_deq_bits_btb_taken),
    .io_deq_bits_btb_bridx(fq_io_deq_bits_btb_bridx),
    .io_deq_bits_btb_entry(fq_io_deq_bits_btb_entry),
    .io_deq_bits_btb_bht_history(fq_io_deq_bits_btb_bht_history),
    .io_deq_bits_pc(fq_io_deq_bits_pc),
    .io_deq_bits_data(fq_io_deq_bits_data),
    .io_deq_bits_xcpt_pf_inst(fq_io_deq_bits_xcpt_pf_inst),
    .io_deq_bits_xcpt_ae_inst(fq_io_deq_bits_xcpt_ae_inst),
    .io_deq_bits_replay(fq_io_deq_bits_replay),
    .io_mask(fq_io_mask),
    .io_covSum(fq_io_covSum),
    .metaAssert(fq_metaAssert),
    .metaReset(fq_metaReset)
  );
  TLB_1 tlb ( // @[Frontend.scala 100:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vaddr(tlb_io_req_bits_vaddr),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_paddr(tlb_io_resp_paddr),
    .io_resp_pf_inst(tlb_io_resp_pf_inst),
    .io_resp_ae_inst(tlb_io_resp_ae_inst),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_sfence_valid(tlb_io_sfence_valid),
    .io_sfence_bits_rs1(tlb_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(tlb_io_sfence_bits_rs2),
    .io_sfence_bits_addr(tlb_io_sfence_bits_addr),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_valid(tlb_io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr(tlb_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(tlb_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(tlb_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(tlb_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(tlb_io_ptw_ptbr_mode),
    .io_ptw_status_debug(tlb_io_ptw_status_debug),
    .io_ptw_status_prv(tlb_io_ptw_status_prv),
    .io_ptw_pmp_0_cfg_l(tlb_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(tlb_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(tlb_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(tlb_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(tlb_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(tlb_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(tlb_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(tlb_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(tlb_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(tlb_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(tlb_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(tlb_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(tlb_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(tlb_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(tlb_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(tlb_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(tlb_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(tlb_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(tlb_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(tlb_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(tlb_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(tlb_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(tlb_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(tlb_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(tlb_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(tlb_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(tlb_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(tlb_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(tlb_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(tlb_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(tlb_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(tlb_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(tlb_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(tlb_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(tlb_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(tlb_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(tlb_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(tlb_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(tlb_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(tlb_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(tlb_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(tlb_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(tlb_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(tlb_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(tlb_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(tlb_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(tlb_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(tlb_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(tlb_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(tlb_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(tlb_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(tlb_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(tlb_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(tlb_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(tlb_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(tlb_io_ptw_pmp_7_mask),
    .io_kill(tlb_io_kill),
    .io_covSum(tlb_io_covSum),
    .metaAssert(tlb_metaAssert),
    .metaReset(tlb_metaReset)
  );
  BTB btb ( // @[Frontend.scala 181:21]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_req_bits_addr(btb_io_req_bits_addr),
    .io_resp_valid(btb_io_resp_valid),
    .io_resp_bits_taken(btb_io_resp_bits_taken),
    .io_resp_bits_bridx(btb_io_resp_bits_bridx),
    .io_resp_bits_target(btb_io_resp_bits_target),
    .io_resp_bits_entry(btb_io_resp_bits_entry),
    .io_resp_bits_bht_history(btb_io_resp_bits_bht_history),
    .io_resp_bits_bht_value(btb_io_resp_bits_bht_value),
    .io_btb_update_valid(btb_io_btb_update_valid),
    .io_btb_update_bits_prediction_entry(btb_io_btb_update_bits_prediction_entry),
    .io_btb_update_bits_pc(btb_io_btb_update_bits_pc),
    .io_btb_update_bits_isValid(btb_io_btb_update_bits_isValid),
    .io_btb_update_bits_br_pc(btb_io_btb_update_bits_br_pc),
    .io_btb_update_bits_cfiType(btb_io_btb_update_bits_cfiType),
    .io_bht_update_valid(btb_io_bht_update_valid),
    .io_bht_update_bits_prediction_history(btb_io_bht_update_bits_prediction_history),
    .io_bht_update_bits_pc(btb_io_bht_update_bits_pc),
    .io_bht_update_bits_branch(btb_io_bht_update_bits_branch),
    .io_bht_update_bits_taken(btb_io_bht_update_bits_taken),
    .io_bht_update_bits_mispredict(btb_io_bht_update_bits_mispredict),
    .io_bht_advance_valid(btb_io_bht_advance_valid),
    .io_bht_advance_bits_bht_value(btb_io_bht_advance_bits_bht_value),
    .io_ras_update_valid(btb_io_ras_update_valid),
    .io_ras_update_bits_cfiType(btb_io_ras_update_bits_cfiType),
    .io_ras_update_bits_returnAddr(btb_io_ras_update_bits_returnAddr),
    .io_ras_head_valid(btb_io_ras_head_valid),
    .io_ras_head_bits(btb_io_ras_head_bits),
    .io_flush(btb_io_flush),
    .io_covSum(btb_io_covSum),
    .metaAssert(btb_metaAssert),
    .metaReset(btb_metaReset)
  );
  assign _T_2 = io_cpu_req_valid | io_cpu_sfence_valid; // @[Frontend.scala 91:29]
  assign _T_3 = _T_2 | io_cpu_flush_icache; // @[Frontend.scala 91:52]
  assign _T_4 = _T_3 | io_cpu_bht_update_valid; // @[Frontend.scala 91:75]
  assign _T_5 = _T_4 | io_cpu_btb_update_valid; // @[Frontend.scala 91:102]
  assign _T_7 = ~_T_5 | io_cpu_might_request; // @[Frontend.scala 91:130]
  assign _T_9 = _T_7 | reset; // @[Frontend.scala 91:9]
  assign _T_17 = ~s1_valid | ~s2_valid; // @[Frontend.scala 106:55]
  assign _T_18 = ~fq_io_mask[3] & _T_17; // @[Frontend.scala 106:41]
  assign _T_19 = ~fq_io_mask[2] | _T_18; // @[Frontend.scala 105:40]
  assign _T_24 = ~s1_valid & ~s2_valid; // @[Frontend.scala 107:55]
  assign _T_25 = ~fq_io_mask[4] & _T_24; // @[Frontend.scala 107:41]
  assign s0_fq_has_space = _T_19 | _T_25; // @[Frontend.scala 106:70]
  assign s0_valid = io_cpu_req_valid | s0_fq_has_space; // @[Frontend.scala 108:35]
  assign _T_27 = ~auto_reset_vector_sink_in | 32'h1; // @[Frontend.scala 343:33]
  assign s2_btb_taken = s2_btb_resp_valid & s2_btb_resp_bits_taken; // @[Frontend.scala 115:40]
  assign s2_xcpt = s2_tlb_resp_ae_inst | s2_tlb_resp_pf_inst; // @[Frontend.scala 117:37]
  assign _T_30 = ~s1_pc | 40'h3; // @[Frontend.scala 123:29]
  assign s1_base_pc = ~_T_30; // @[Frontend.scala 123:20]
  assign ntpc = s1_base_pc + 40'h4; // @[Frontend.scala 124:25]
  assign _T_32 = fq_io_enq_ready & fq_io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_34 = s2_valid & ~_T_32; // @[Frontend.scala 129:26]
  assign s2_replay = _T_34 | _T_37; // @[Frontend.scala 129:48]
  assign _T_36 = s2_replay & ~s0_valid; // @[Frontend.scala 129:69]
  assign _T_105 = s2_partial_insn[1:0] != 2'h3; // @[Frontend.scala 210:45]
  assign taken_prevRVI = s2_partial_insn_valid & ~_T_105; // @[Frontend.scala 211:31]
  assign taken_bits = fq_io_enq_bits_data[15:0]; // @[Frontend.scala 213:37]
  assign taken_rviBits = {taken_bits,s2_partial_insn}; // @[Cat.scala 29:58]
  assign taken_rviJump = taken_rviBits[6:0] == 7'h6f; // @[Frontend.scala 217:34]
  assign taken_rviJALR = taken_rviBits[6:0] == 7'h67; // @[Frontend.scala 218:34]
  assign _T_299 = taken_rviJump | taken_rviJALR; // @[Frontend.scala 232:29]
  assign taken_rviBranch = taken_rviBits[6:0] == 7'h63; // @[Frontend.scala 216:36]
  assign _T_300 = taken_rviBranch & s2_btb_resp_bits_bht_value; // @[Frontend.scala 232:53]
  assign _T_301 = _T_299 | _T_300; // @[Frontend.scala 232:40]
  assign _T_302 = taken_prevRVI & _T_301; // @[Frontend.scala 232:17]
  assign taken_valid = fq_io_enq_bits_mask[0] & ~taken_prevRVI; // @[Frontend.scala 212:44]
  assign _T_127 = taken_bits & 16'he003; // @[Frontend.scala 223:26]
  assign taken_rvcJump = 16'ha001 == _T_127; // @[Frontend.scala 223:26]
  assign _T_169 = taken_bits & 16'hf003; // @[Frontend.scala 227:26]
  assign _T_170 = 16'h9002 == _T_169; // @[Frontend.scala 227:26]
  assign _T_172 = taken_bits[6:2] == 5'h0; // @[Frontend.scala 227:62]
  assign taken_rvcJALR = _T_170 & _T_172; // @[Frontend.scala 227:49]
  assign _T_303 = taken_rvcJump | taken_rvcJALR; // @[Frontend.scala 233:27]
  assign _T_163 = 16'h8002 == _T_169; // @[Frontend.scala 225:24]
  assign taken_rvcJR = _T_163 & _T_172; // @[Frontend.scala 225:46]
  assign _T_304 = _T_303 | taken_rvcJR; // @[Frontend.scala 233:38]
  assign _T_122 = 16'hc001 == _T_127; // @[Frontend.scala 221:28]
  assign _T_124 = 16'he001 == _T_127; // @[Frontend.scala 221:60]
  assign taken_rvcBranch = _T_122 | _T_124; // @[Frontend.scala 221:52]
  assign _T_305 = taken_rvcBranch & s2_btb_resp_bits_bht_value; // @[Frontend.scala 233:60]
  assign _T_306 = _T_304 | _T_305; // @[Frontend.scala 233:47]
  assign _T_307 = taken_valid & _T_306; // @[Frontend.scala 233:15]
  assign taken_taken = _T_302 | _T_307; // @[Frontend.scala 232:71]
  assign taken_idx = ~taken_taken; // @[Frontend.scala 247:13]
  assign _T_372 = taken_bits[1:0] != 2'h3; // @[Frontend.scala 210:45]
  assign taken_prevRVI_1 = taken_valid & ~_T_372; // @[Frontend.scala 211:31]
  assign taken_bits_1 = fq_io_enq_bits_data[31:16]; // @[Frontend.scala 213:37]
  assign taken_rviBits_1 = {taken_bits_1,taken_bits}; // @[Cat.scala 29:58]
  assign taken_rviJALR_1 = taken_rviBits_1[6:0] == 7'h67; // @[Frontend.scala 218:34]
  assign _T_382 = taken_rviJALR_1 & ~taken_rviBits_1[7]; // @[Frontend.scala 219:31]
  assign _T_384 = taken_rviBits_1[19:15] & 5'h1b; // @[Frontend.scala 219:66]
  assign _T_385 = 5'h1 == _T_384; // @[Frontend.scala 219:66]
  assign taken_rviReturn_1 = _T_382 & _T_385; // @[Frontend.scala 219:46]
  assign _T_575 = taken_prevRVI_1 & taken_rviReturn_1; // @[Frontend.scala 234:61]
  assign taken_valid_1 = fq_io_enq_bits_mask[1] & ~taken_prevRVI_1; // @[Frontend.scala 212:44]
  assign _T_429 = taken_bits_1 & 16'hf003; // @[Frontend.scala 225:24]
  assign _T_430 = 16'h8002 == _T_429; // @[Frontend.scala 225:24]
  assign _T_432 = taken_bits_1[6:2] == 5'h0; // @[Frontend.scala 225:59]
  assign taken_rvcJR_1 = _T_430 & _T_432; // @[Frontend.scala 225:46]
  assign _T_434 = taken_bits_1[11:7] & 5'h1b; // @[Frontend.scala 226:49]
  assign _T_435 = 5'h1 == _T_434; // @[Frontend.scala 226:49]
  assign taken_rvcReturn_1 = taken_rvcJR_1 & _T_435; // @[Frontend.scala 226:29]
  assign _T_576 = taken_valid_1 & taken_rvcReturn_1; // @[Frontend.scala 234:83]
  assign _T_577 = _T_575 | _T_576; // @[Frontend.scala 234:74]
  assign taken_predictReturn_1 = btb_io_ras_head_valid & _T_577; // @[Frontend.scala 234:49]
  assign _T_616 = s2_valid & taken_predictReturn_1; // @[Frontend.scala 260:26]
  assign _T_115 = taken_rviJALR & ~taken_rviBits[7]; // @[Frontend.scala 219:31]
  assign _T_117 = taken_rviBits[19:15] & 5'h1b; // @[Frontend.scala 219:66]
  assign _T_118 = 5'h1 == _T_117; // @[Frontend.scala 219:66]
  assign taken_rviReturn = _T_115 & _T_118; // @[Frontend.scala 219:46]
  assign _T_308 = taken_prevRVI & taken_rviReturn; // @[Frontend.scala 234:61]
  assign _T_167 = taken_bits[11:7] & 5'h1b; // @[Frontend.scala 226:49]
  assign _T_168 = 5'h1 == _T_167; // @[Frontend.scala 226:49]
  assign taken_rvcReturn = taken_rvcJR & _T_168; // @[Frontend.scala 226:29]
  assign _T_309 = taken_valid & taken_rvcReturn; // @[Frontend.scala 234:83]
  assign _T_310 = _T_308 | _T_309; // @[Frontend.scala 234:74]
  assign taken_predictReturn = btb_io_ras_head_valid & _T_310; // @[Frontend.scala 234:49]
  assign _T_349 = s2_valid & taken_predictReturn; // @[Frontend.scala 260:26]
  assign _GEN_45 = ~s2_btb_taken & _T_349; // @[Frontend.scala 256:30]
  assign _GEN_78 = _T_616 | _GEN_45; // @[Frontend.scala 260:44]
  assign _GEN_81 = s2_btb_taken ? _GEN_45 : _GEN_78; // @[Frontend.scala 256:30]
  assign useRAS = taken_idx ? _GEN_81 : _GEN_45; // @[Frontend.scala 247:25]
  assign taken_rviBranch_1 = taken_rviBits_1[6:0] == 7'h63; // @[Frontend.scala 216:36]
  assign _T_580 = taken_prevRVI_1 & taken_rviBranch_1; // @[Frontend.scala 236:53]
  assign _T_388 = taken_bits_1 & 16'he003; // @[Frontend.scala 221:28]
  assign _T_389 = 16'hc001 == _T_388; // @[Frontend.scala 221:28]
  assign _T_391 = 16'he001 == _T_388; // @[Frontend.scala 221:60]
  assign taken_rvcBranch_1 = _T_389 | _T_391; // @[Frontend.scala 221:52]
  assign _T_581 = taken_valid_1 & taken_rvcBranch_1; // @[Frontend.scala 236:75]
  assign _T_582 = _T_580 | _T_581; // @[Frontend.scala 236:66]
  assign taken_predictBranch_1 = s2_btb_resp_bits_bht_value & _T_582; // @[Frontend.scala 236:41]
  assign taken_rviJump_1 = taken_rviBits_1[6:0] == 7'h6f; // @[Frontend.scala 217:34]
  assign _T_578 = taken_prevRVI_1 & taken_rviJump_1; // @[Frontend.scala 235:33]
  assign taken_rvcJump_1 = 16'ha001 == _T_388; // @[Frontend.scala 223:26]
  assign _T_579 = taken_valid_1 & taken_rvcJump_1; // @[Frontend.scala 235:53]
  assign taken_predictJump_1 = _T_578 | _T_579; // @[Frontend.scala 235:44]
  assign _T_617 = taken_predictBranch_1 | taken_predictJump_1; // @[Frontend.scala 263:44]
  assign _T_618 = s2_valid & _T_617; // @[Frontend.scala 263:26]
  assign _T_91 = ~s2_pc | 40'h3; // @[Frontend.scala 203:31]
  assign s2_base_pc = ~_T_91; // @[Frontend.scala 203:22]
  assign taken_pc_1 = s2_base_pc | 40'h2; // @[Frontend.scala 264:33]
  assign _T_620 = taken_pc_1 - 40'h2; // @[Frontend.scala 267:36]
  assign _T_622 = taken_prevRVI_1 ? _T_620 : taken_pc_1; // @[Frontend.scala 267:57]
  assign _T_443 = taken_rviBits_1[31]; // @[RocketCore.scala 1036:53]
  assign _T_498 = taken_rviBits_1[31]; // @[Cat.scala 29:58]
  assign _T_497 = {11{_T_443}}; // @[Cat.scala 29:58]
  assign _T_495 = taken_rviBits_1[19:12]; // @[Cat.scala 29:58]
  assign _T_494 = taken_rviBits_1[20]; // @[Cat.scala 29:58]
  assign _T_502 = {_T_498,_T_497,_T_495,_T_494,taken_rviBits_1[30:25],taken_rviBits_1[24:21],1'h0}; // @[RocketCore.scala 1050:53]
  assign _T_557 = {8{_T_443}}; // @[Cat.scala 29:58]
  assign _T_556 = taken_rviBits_1[7]; // @[Cat.scala 29:58]
  assign _T_564 = {_T_498,_T_497,_T_557,_T_556,taken_rviBits_1[30:25],taken_rviBits_1[11:8],1'h0}; // @[RocketCore.scala 1050:53]
  assign taken_rviImm_1 = taken_rviBits_1[3] ? $signed(_T_502) : $signed(_T_564); // @[Frontend.scala 229:23]
  assign _T_399 = taken_bits_1[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  assign _T_409 = {_T_399,taken_bits_1[6:5],taken_bits_1[2],taken_bits_1[11:10],taken_bits_1[4:3],1'h0}; // @[Frontend.scala 224:66]
  assign _T_412 = taken_bits_1[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  assign _T_428 = {_T_412,taken_bits_1[8],taken_bits_1[10:9],taken_bits_1[6],taken_bits_1[7],taken_bits_1[2],taken_bits_1[11],taken_bits_1[5:3],1'h0}; // @[Frontend.scala 224:106]
  assign taken_rvcImm_1 = taken_bits_1[14] ? $signed({{8{_T_409[12]}},_T_409}) : $signed(_T_428); // @[Frontend.scala 224:23]
  assign _T_623 = taken_prevRVI_1 ? $signed(taken_rviImm_1) : $signed({{11{taken_rvcImm_1[20]}},taken_rvcImm_1}); // @[Frontend.scala 267:69]
  assign _GEN_127 = {{8{_T_623[31]}},_T_623}; // @[Frontend.scala 267:64]
  assign _T_626 = $signed(_T_622) + $signed(_GEN_127); // @[Frontend.scala 268:34]
  assign _T_313 = taken_prevRVI & taken_rviBranch; // @[Frontend.scala 236:53]
  assign _T_314 = taken_valid & taken_rvcBranch; // @[Frontend.scala 236:75]
  assign _T_315 = _T_313 | _T_314; // @[Frontend.scala 236:66]
  assign taken_predictBranch = s2_btb_resp_bits_bht_value & _T_315; // @[Frontend.scala 236:41]
  assign _T_311 = taken_prevRVI & taken_rviJump; // @[Frontend.scala 235:33]
  assign _T_312 = taken_valid & taken_rvcJump; // @[Frontend.scala 235:53]
  assign taken_predictJump = _T_311 | _T_312; // @[Frontend.scala 235:44]
  assign _T_350 = taken_predictBranch | taken_predictJump; // @[Frontend.scala 263:44]
  assign _T_351 = s2_valid & _T_350; // @[Frontend.scala 263:26]
  assign _T_352 = ~_T_91; // @[Frontend.scala 266:32]
  assign _T_176 = taken_rviBits[31]; // @[RocketCore.scala 1036:53]
  assign _T_231 = taken_rviBits[31]; // @[Cat.scala 29:58]
  assign _T_230 = {11{_T_176}}; // @[Cat.scala 29:58]
  assign _T_228 = taken_rviBits[19:12]; // @[Cat.scala 29:58]
  assign _T_227 = taken_rviBits[20]; // @[Cat.scala 29:58]
  assign _T_235 = {_T_231,_T_230,_T_228,_T_227,taken_rviBits[30:25],taken_rviBits[24:21],1'h0}; // @[RocketCore.scala 1050:53]
  assign _T_290 = {8{_T_176}}; // @[Cat.scala 29:58]
  assign _T_289 = taken_rviBits[7]; // @[Cat.scala 29:58]
  assign _T_297 = {_T_231,_T_230,_T_290,_T_289,taken_rviBits[30:25],taken_rviBits[11:8],1'h0}; // @[RocketCore.scala 1050:53]
  assign taken_rviImm = taken_rviBits[3] ? $signed(_T_235) : $signed(_T_297); // @[Frontend.scala 229:23]
  assign _T_353 = $signed(taken_rviImm) - 32'sh2; // @[Frontend.scala 266:61]
  assign _T_132 = taken_bits[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  assign _T_142 = {_T_132,taken_bits[6:5],taken_bits[2],taken_bits[11:10],taken_bits[4:3],1'h0}; // @[Frontend.scala 224:66]
  assign _T_145 = taken_bits[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  assign _T_161 = {_T_145,taken_bits[8],taken_bits[10:9],taken_bits[6],taken_bits[7],taken_bits[2],taken_bits[11],taken_bits[5:3],1'h0}; // @[Frontend.scala 224:106]
  assign taken_rvcImm = taken_bits[14] ? $signed({{8{_T_142[12]}},_T_142}) : $signed(_T_161); // @[Frontend.scala 224:23]
  assign _T_354 = taken_prevRVI ? $signed(_T_353) : $signed({{12{taken_rvcImm[20]}},taken_rvcImm}); // @[Frontend.scala 266:44]
  assign _GEN_128 = {{7{_T_354[32]}},_T_354}; // @[Frontend.scala 266:39]
  assign _T_357 = $signed(_T_352) + $signed(_GEN_128); // @[Frontend.scala 268:34]
  assign predicted_taken = btb_io_resp_valid & btb_io_resp_bits_taken; // @[Frontend.scala 194:29]
  assign _T_89 = {btb_io_resp_bits_target[38],btb_io_resp_bits_target}; // @[Cat.scala 29:58]
  assign _GEN_28 = predicted_taken ? _T_89 : ntpc; // @[Frontend.scala 194:56]
  assign _GEN_43 = _T_351 ? _T_357 : _GEN_28; // @[Frontend.scala 263:61]
  assign _GEN_46 = s2_btb_taken ? _GEN_28 : _GEN_43; // @[Frontend.scala 256:30]
  assign _GEN_79 = _T_618 ? _T_626 : _GEN_46; // @[Frontend.scala 263:61]
  assign _GEN_82 = s2_btb_taken ? _GEN_46 : _GEN_79; // @[Frontend.scala 256:30]
  assign _GEN_99 = taken_idx ? _GEN_82 : _GEN_46; // @[Frontend.scala 247:25]
  assign predicted_npc = useRAS ? {{1'd0}, btb_io_ras_head_bits} : _GEN_99; // @[Frontend.scala 307:19]
  assign npc = s2_replay ? s2_pc : predicted_npc; // @[Frontend.scala 130:16]
  assign _T_40 = s2_valid & ~s2_speculative; // @[Frontend.scala 136:53]
  assign _T_41 = s1_speculative | _T_40; // @[Frontend.scala 136:41]
  assign s0_speculative = _T_41 | predicted_taken; // @[Frontend.scala 136:72]
  assign _T_566 = taken_rviJump_1 | taken_rviJALR_1; // @[Frontend.scala 232:29]
  assign _T_567 = taken_rviBranch_1 & s2_btb_resp_bits_bht_value; // @[Frontend.scala 232:53]
  assign _T_568 = _T_566 | _T_567; // @[Frontend.scala 232:40]
  assign _T_569 = taken_prevRVI_1 & _T_568; // @[Frontend.scala 232:17]
  assign _T_437 = 16'h9002 == _T_429; // @[Frontend.scala 227:26]
  assign taken_rvcJALR_1 = _T_437 & _T_432; // @[Frontend.scala 227:49]
  assign _T_570 = taken_rvcJump_1 | taken_rvcJALR_1; // @[Frontend.scala 233:27]
  assign _T_571 = _T_570 | taken_rvcJR_1; // @[Frontend.scala 233:38]
  assign _T_572 = taken_rvcBranch_1 & s2_btb_resp_bits_bht_value; // @[Frontend.scala 233:60]
  assign _T_573 = _T_571 | _T_572; // @[Frontend.scala 233:47]
  assign _T_574 = taken_valid_1 & _T_573; // @[Frontend.scala 233:15]
  assign taken_taken_1 = _T_569 | _T_574; // @[Frontend.scala 232:71]
  assign taken = taken_taken | taken_taken_1; // @[Frontend.scala 288:19]
  assign _GEN_116 = _T_32 | io_cpu_req_valid; // @[Frontend.scala 318:33]
  assign _GEN_120 = taken ? _GEN_116 : io_cpu_req_valid; // @[Frontend.scala 314:20]
  assign s2_redirect = s2_btb_taken ? io_cpu_req_valid : _GEN_120; // @[Frontend.scala 313:26]
  assign _GEN_0 = ~s2_replay & ~s2_redirect; // @[Frontend.scala 142:21]
  assign _T_49 = s2_redirect | tlb_io_resp_miss; // @[Frontend.scala 162:36]
  assign s2_can_speculatively_refill = s2_tlb_resp_cacheable & ~io_ptw_customCSRs_csrs_0_value[3]; // @[Frontend.scala 163:59]
  assign _T_54 = s2_speculative & ~s2_can_speculatively_refill; // @[Frontend.scala 164:39]
  assign _T_60 = _T_59 & s2_valid; // @[Frontend.scala 167:40]
  assign _T_62 = ~s2_tlb_resp_miss & icache_io_s2_kill; // @[Frontend.scala 167:98]
  assign _T_63 = icache_io_resp_valid | _T_62; // @[Frontend.scala 167:77]
  assign _T_65 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc; // @[Frontend.scala 169:28]
  assign _T_67 = ~_T_65 | 40'h1; // @[Frontend.scala 343:33]
  assign _T_70 = 3'h3 << s2_pc[1]; // @[Frontend.scala 172:52]
  assign _T_72 = icache_io_s2_kill & ~icache_io_resp_valid; // @[Frontend.scala 173:76]
  assign _T_74 = _T_72 & ~s2_xcpt; // @[Frontend.scala 173:101]
  assign _T_75 = icache_io_resp_bits_replay | _T_74; // @[Frontend.scala 173:55]
  assign _T_77 = s2_speculative & io_ptw_customCSRs_csrs_0_value[3]; // @[Frontend.scala 177:27]
  assign _T_79 = _T_77 & ~icache_io_s2_kill; // @[Frontend.scala 177:110]
  assign _T_82 = ~_T_79 | reset; // @[Frontend.scala 177:9]
  assign _T_84 = icache_io_resp_valid & icache_io_resp_bits_ae; // @[Frontend.scala 178:30]
  assign fetch_bubble_likely = ~fq_io_mask[1]; // @[Frontend.scala 295:33]
  assign _T_96 = _T_32 & ~wrong_path; // @[Frontend.scala 296:51]
  assign _T_97 = _T_96 & fetch_bubble_likely; // @[Frontend.scala 296:66]
  assign _T_635 = taken_predictBranch_1 & s2_btb_resp_bits_bht_value; // @[Frontend.scala 275:52]
  assign _T_636 = _T_635 | taken_predictJump_1; // @[Frontend.scala 275:91]
  assign _T_637 = _T_636 | taken_predictReturn_1; // @[Frontend.scala 275:106]
  assign _T_638 = ~s2_btb_resp_valid & _T_637; // @[Frontend.scala 275:34]
  assign _T_366 = taken_predictBranch & s2_btb_resp_bits_bht_value; // @[Frontend.scala 275:52]
  assign _T_367 = _T_366 | taken_predictJump; // @[Frontend.scala 275:91]
  assign _T_368 = _T_367 | taken_predictReturn; // @[Frontend.scala 275:106]
  assign _T_369 = ~s2_btb_resp_valid & _T_368; // @[Frontend.scala 275:34]
  assign _GEN_92 = _T_638 | _T_369; // @[Frontend.scala 275:125]
  assign updateBTB = taken_idx ? _GEN_92 : _T_369; // @[Frontend.scala 247:25]
  assign _T_98 = _T_97 & updateBTB; // @[Frontend.scala 296:89]
  assign _T_99 = {taken_idx, 1'h0}; // @[Frontend.scala 300:63]
  assign _GEN_129 = {{38'd0}, _T_99}; // @[Frontend.scala 300:50]
  assign _T_100 = s2_base_pc | _GEN_129; // @[Frontend.scala 300:50]
  assign _GEN_36 = io_cpu_btb_update_valid ? {{1'd0}, io_cpu_btb_update_bits_br_pc} : _T_100; // @[Frontend.scala 294:37]
  assign _GEN_37 = io_cpu_btb_update_valid ? {{1'd0}, io_cpu_btb_update_bits_pc} : s2_base_pc; // @[Frontend.scala 294:37]
  assign after_idx = taken_idx ? 2'h2 : 2'h1; // @[Frontend.scala 247:25]
  assign _T_101 = {after_idx, 1'h0}; // @[Frontend.scala 304:66]
  assign _GEN_130 = {{37'd0}, _T_101}; // @[Frontend.scala 304:53]
  assign _T_103 = s2_base_pc + _GEN_130; // @[Frontend.scala 304:53]
  assign _T_119 = taken_rviJALR | taken_rviJump; // @[Frontend.scala 220:30]
  assign taken_rviCall = _T_119 & taken_rviBits[7]; // @[Frontend.scala 220:42]
  assign _T_316 = s2_valid & s2_btb_resp_valid; // @[Frontend.scala 238:22]
  assign _T_318 = _T_316 & ~s2_btb_resp_bits_bridx; // @[Frontend.scala 238:43]
  assign _T_319 = _T_318 & taken_valid; // @[Frontend.scala 238:77]
  assign _T_321 = _T_319 & ~_T_372; // @[Frontend.scala 238:86]
  assign _GEN_39 = _T_321 | _T_75; // @[Frontend.scala 238:95]
  assign _GEN_40 = _T_321 | wrong_path; // @[Frontend.scala 238:95]
  assign _T_326 = taken_rviCall | taken_rviReturn; // @[Frontend.scala 250:92]
  assign _T_327 = taken_prevRVI & _T_326; // @[Frontend.scala 250:80]
  assign _T_328 = taken_rvcJALR | taken_rvcReturn; // @[Frontend.scala 250:127]
  assign _T_329 = taken_valid & _T_328; // @[Frontend.scala 250:115]
  assign _T_330 = _T_327 | _T_329; // @[Frontend.scala 250:106]
  assign _T_331 = _T_96 & _T_330; // @[Frontend.scala 250:68]
  assign _T_332 = taken_prevRVI ? taken_rviReturn : taken_rvcReturn; // @[Frontend.scala 251:50]
  assign _T_333 = taken_prevRVI ? taken_rviCall : taken_rvcJALR; // @[Frontend.scala 252:50]
  assign _T_334 = taken_prevRVI ? taken_rviBranch : taken_rvcBranch; // @[Frontend.scala 253:50]
  assign _T_337 = _T_334 ? 1'h0 : 1'h1; // @[Frontend.scala 253:46]
  assign _T_338 = _T_333 ? 2'h2 : {{1'd0}, _T_337}; // @[Frontend.scala 252:46]
  assign _T_339 = _T_332 ? 2'h3 : _T_338; // @[Frontend.scala 251:46]
  assign _T_342 = _T_32 & taken_taken; // @[Frontend.scala 257:34]
  assign _T_344 = _T_342 & ~taken_predictBranch; // @[Frontend.scala 257:43]
  assign _T_346 = _T_344 & ~taken_predictJump; // @[Frontend.scala 257:61]
  assign _T_348 = _T_346 & ~taken_predictReturn; // @[Frontend.scala 257:77]
  assign _GEN_41 = _T_348 | _GEN_40; // @[Frontend.scala 257:96]
  assign _GEN_44 = s2_btb_taken ? _GEN_40 : _GEN_41; // @[Frontend.scala 256:30]
  assign _GEN_47 = _T_315 & _T_96; // @[Frontend.scala 271:59]
  assign taken_rvc_1 = taken_bits_1[1:0] != 2'h3; // @[Frontend.scala 210:45]
  assign _T_386 = taken_rviJALR_1 | taken_rviJump_1; // @[Frontend.scala 220:30]
  assign taken_rviCall_1 = _T_386 & taken_rviBits_1[7]; // @[Frontend.scala 220:42]
  assign _T_585 = _T_316 & s2_btb_resp_bits_bridx; // @[Frontend.scala 238:43]
  assign _T_586 = _T_585 & taken_valid_1; // @[Frontend.scala 238:77]
  assign _T_588 = _T_586 & ~taken_rvc_1; // @[Frontend.scala 238:86]
  assign _GEN_76 = _T_588 | _GEN_44; // @[Frontend.scala 238:95]
  assign _T_593 = taken_rviCall_1 | taken_rviReturn_1; // @[Frontend.scala 250:92]
  assign _T_594 = taken_prevRVI_1 & _T_593; // @[Frontend.scala 250:80]
  assign _T_595 = taken_rvcJALR_1 | taken_rvcReturn_1; // @[Frontend.scala 250:127]
  assign _T_596 = taken_valid_1 & _T_595; // @[Frontend.scala 250:115]
  assign _T_597 = _T_594 | _T_596; // @[Frontend.scala 250:106]
  assign _T_598 = _T_96 & _T_597; // @[Frontend.scala 250:68]
  assign _T_599 = taken_prevRVI_1 ? taken_rviReturn_1 : taken_rvcReturn_1; // @[Frontend.scala 251:50]
  assign _T_600 = taken_prevRVI_1 ? taken_rviCall_1 : taken_rvcJALR_1; // @[Frontend.scala 252:50]
  assign _T_601 = taken_prevRVI_1 ? taken_rviBranch_1 : taken_rvcBranch_1; // @[Frontend.scala 253:50]
  assign _T_604 = _T_601 ? 1'h0 : 1'h1; // @[Frontend.scala 253:46]
  assign _T_605 = _T_600 ? 2'h2 : {{1'd0}, _T_604}; // @[Frontend.scala 252:46]
  assign _T_606 = _T_599 ? 2'h3 : _T_605; // @[Frontend.scala 251:46]
  assign _T_609 = _T_32 & taken_taken_1; // @[Frontend.scala 257:34]
  assign _T_611 = _T_609 & ~taken_predictBranch_1; // @[Frontend.scala 257:43]
  assign _T_613 = _T_611 & ~taken_predictJump_1; // @[Frontend.scala 257:61]
  assign _T_615 = _T_613 & ~taken_predictReturn_1; // @[Frontend.scala 257:77]
  assign _GEN_77 = _T_615 | _GEN_76; // @[Frontend.scala 257:96]
  assign _GEN_83 = _T_582 ? _T_96 : _GEN_47; // @[Frontend.scala 271:59]
  assign _T_641 = taken_valid_1 & taken_idx; // @[Frontend.scala 283:23]
  assign _T_643 = _T_641 & ~taken_rvc_1; // @[Frontend.scala 283:37]
  assign _T_644 = taken_bits_1 | 16'h3; // @[Frontend.scala 285:37]
  assign _T_646 = s2_btb_taken | taken; // @[Frontend.scala 310:45]
  assign _T_647 = _T_32 & _T_646; // @[Frontend.scala 310:28]
  assign _GEN_117 = taken ? taken_idx : s2_btb_resp_bits_bridx; // @[Frontend.scala 314:20]
  assign _GEN_118 = taken | s2_btb_taken; // @[Frontend.scala 314:20]
  assign _GEN_119 = taken ? 5'h1c : s2_btb_resp_bits_entry; // @[Frontend.scala 314:20]
  assign _T_652 = ~s2_partial_insn_valid | fq_io_enq_bits_mask[0]; // @[Frontend.scala 322:35]
  assign _T_654 = _T_652 | reset; // @[Frontend.scala 322:11]
  assign auto_icache_master_out_a_valid = icache_auto_master_out_a_valid; // @[LazyModule.scala 305:12]
  assign auto_icache_master_out_a_bits_address = icache_auto_master_out_a_bits_address; // @[LazyModule.scala 305:12]
  assign io_cpu_resp_valid = fq_io_deq_valid; // @[Frontend.scala 327:15]
  assign io_cpu_resp_bits_btb_taken = fq_io_deq_bits_btb_taken; // @[Frontend.scala 327:15]
  assign io_cpu_resp_bits_btb_bridx = fq_io_deq_bits_btb_bridx; // @[Frontend.scala 327:15]
  assign io_cpu_resp_bits_btb_entry = fq_io_deq_bits_btb_entry; // @[Frontend.scala 327:15]
  assign io_cpu_resp_bits_btb_bht_history = fq_io_deq_bits_btb_bht_history; // @[Frontend.scala 327:15]
  assign io_cpu_resp_bits_pc = fq_io_deq_bits_pc; // @[Frontend.scala 327:15]
  assign io_cpu_resp_bits_data = fq_io_deq_bits_data; // @[Frontend.scala 327:15]
  assign io_cpu_resp_bits_xcpt_pf_inst = fq_io_deq_bits_xcpt_pf_inst; // @[Frontend.scala 327:15]
  assign io_cpu_resp_bits_xcpt_ae_inst = fq_io_deq_bits_xcpt_ae_inst; // @[Frontend.scala 327:15]
  assign io_cpu_resp_bits_replay = fq_io_deq_bits_replay; // @[Frontend.scala 327:15]
  assign io_cpu_npc = ~_T_67; // @[Frontend.scala 169:14]
  assign io_ptw_req_valid = tlb_io_ptw_req_valid; // @[Frontend.scala 149:10]
  assign io_ptw_req_bits_valid = tlb_io_ptw_req_bits_valid; // @[Frontend.scala 149:10]
  assign io_ptw_req_bits_bits_addr = tlb_io_ptw_req_bits_bits_addr; // @[Frontend.scala 149:10]
  assign icache_clock = gated_clock; // @[Frontend.scala 96:16]
  assign icache_reset = reset;
  assign icache_auto_master_out_a_ready = auto_icache_master_out_a_ready; // @[LazyModule.scala 305:12]
  assign icache_auto_master_out_d_valid = auto_icache_master_out_d_valid; // @[LazyModule.scala 305:12]
  assign icache_auto_master_out_d_bits_opcode = auto_icache_master_out_d_bits_opcode; // @[LazyModule.scala 305:12]
  assign icache_auto_master_out_d_bits_size = auto_icache_master_out_d_bits_size; // @[LazyModule.scala 305:12]
  assign icache_auto_master_out_d_bits_data = auto_icache_master_out_d_bits_data; // @[LazyModule.scala 305:12]
  assign icache_auto_master_out_d_bits_corrupt = auto_icache_master_out_d_bits_corrupt; // @[LazyModule.scala 305:12]
  assign icache_io_req_valid = io_cpu_req_valid | s0_fq_has_space; // @[Frontend.scala 157:23]
  assign icache_io_req_bits_addr = io_cpu_npc[38:0]; // @[Frontend.scala 158:27]
  assign icache_io_s1_paddr = tlb_io_resp_paddr; // @[Frontend.scala 160:22]
  assign icache_io_s1_kill = _T_49 | s2_replay; // @[Frontend.scala 162:21]
  assign icache_io_s2_kill = _T_54 | s2_xcpt; // @[Frontend.scala 164:21]
  assign icache_io_invalidate = io_cpu_flush_icache; // @[Frontend.scala 159:24]
  assign fq_clock = gated_clock;
  assign fq_reset = reset | io_cpu_req_valid;
  assign fq_io_enq_valid = _T_60 & _T_63; // @[Frontend.scala 167:19]
  assign fq_io_enq_bits_btb_taken = s2_btb_taken ? s2_btb_taken : _GEN_118; // @[Frontend.scala 174:22 Frontend.scala 175:28 Frontend.scala 316:34]
  assign fq_io_enq_bits_btb_bridx = s2_btb_taken ? s2_btb_resp_bits_bridx : _GEN_117; // @[Frontend.scala 174:22 Frontend.scala 315:34]
  assign fq_io_enq_bits_btb_entry = s2_btb_taken ? s2_btb_resp_bits_entry : _GEN_119; // @[Frontend.scala 174:22 Frontend.scala 317:34]
  assign fq_io_enq_bits_btb_bht_history = s2_btb_resp_bits_bht_history; // @[Frontend.scala 174:22]
  assign fq_io_enq_bits_pc = s2_pc; // @[Frontend.scala 168:21]
  assign fq_io_enq_bits_data = icache_io_resp_bits_data; // @[Frontend.scala 171:23]
  assign fq_io_enq_bits_mask = _T_70[1:0]; // @[Frontend.scala 172:23]
  assign fq_io_enq_bits_xcpt_pf_inst = s2_tlb_resp_pf_inst; // @[Frontend.scala 176:23]
  assign fq_io_enq_bits_xcpt_ae_inst = _T_84 | s2_tlb_resp_ae_inst; // @[Frontend.scala 176:23 Frontend.scala 178:87]
  assign fq_io_enq_bits_replay = _T_588 | _GEN_39; // @[Frontend.scala 173:25 Frontend.scala 242:31 Frontend.scala 242:31]
  assign fq_io_deq_ready = io_cpu_resp_ready; // @[Frontend.scala 327:15]
  assign tlb_clock = gated_clock;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = s1_valid & ~s2_replay; // @[Frontend.scala 150:20]
  assign tlb_io_req_bits_vaddr = s1_pc; // @[Frontend.scala 151:25]
  assign tlb_io_sfence_valid = io_cpu_sfence_valid; // @[Frontend.scala 154:17]
  assign tlb_io_sfence_bits_rs1 = io_cpu_sfence_bits_rs1; // @[Frontend.scala 154:17]
  assign tlb_io_sfence_bits_rs2 = io_cpu_sfence_bits_rs2; // @[Frontend.scala 154:17]
  assign tlb_io_sfence_bits_addr = io_cpu_sfence_bits_addr; // @[Frontend.scala 154:17]
  assign tlb_io_ptw_req_ready = io_ptw_req_ready; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_bits_ae = io_ptw_resp_bits_ae; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_bits_level = io_ptw_resp_bits_level; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_resp_bits_homogeneous = io_ptw_resp_bits_homogeneous; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_ptbr_mode = io_ptw_ptbr_mode; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_status_debug = io_ptw_status_debug; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_status_prv = io_ptw_status_prv; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr; // @[Frontend.scala 149:10]
  assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask; // @[Frontend.scala 149:10]
  assign tlb_io_kill = ~s2_valid; // @[Frontend.scala 155:15]
  assign btb_clock = gated_clock;
  assign btb_reset = reset;
  assign btb_io_req_bits_addr = s1_pc[38:0]; // @[Frontend.scala 184:26]
  assign btb_io_btb_update_valid = io_cpu_btb_update_valid ? io_cpu_btb_update_valid : _T_98; // @[Frontend.scala 185:23 Frontend.scala 296:31]
  assign btb_io_btb_update_bits_prediction_entry = io_cpu_btb_update_valid ? io_cpu_btb_update_bits_prediction_entry : 5'h1c; // @[Frontend.scala 185:23 Frontend.scala 297:47]
  assign btb_io_btb_update_bits_pc = _GEN_37[38:0]; // @[Frontend.scala 185:23 Frontend.scala 301:33]
  assign btb_io_btb_update_bits_isValid = ~io_cpu_btb_update_valid | io_cpu_btb_update_bits_isValid; // @[Frontend.scala 185:23 Frontend.scala 298:38]
  assign btb_io_btb_update_bits_br_pc = _GEN_36[38:0]; // @[Frontend.scala 185:23 Frontend.scala 300:36]
  assign btb_io_btb_update_bits_cfiType = io_cpu_btb_update_valid ? io_cpu_btb_update_bits_cfiType : btb_io_ras_update_bits_cfiType; // @[Frontend.scala 185:23 Frontend.scala 299:38]
  assign btb_io_bht_update_valid = io_cpu_bht_update_valid; // @[Frontend.scala 186:23 Frontend.scala 201:50]
  assign btb_io_bht_update_bits_prediction_history = io_cpu_bht_update_bits_prediction_history; // @[Frontend.scala 186:23]
  assign btb_io_bht_update_bits_pc = io_cpu_bht_update_bits_pc; // @[Frontend.scala 186:23]
  assign btb_io_bht_update_bits_branch = io_cpu_bht_update_bits_branch; // @[Frontend.scala 186:23]
  assign btb_io_bht_update_bits_taken = io_cpu_bht_update_bits_taken; // @[Frontend.scala 186:23]
  assign btb_io_bht_update_bits_mispredict = io_cpu_bht_update_bits_mispredict; // @[Frontend.scala 186:23]
  assign btb_io_bht_advance_valid = taken_idx ? _GEN_83 : _GEN_47; // @[Frontend.scala 188:30 Frontend.scala 272:36 Frontend.scala 272:36]
  assign btb_io_bht_advance_bits_bht_value = s2_btb_resp_bits_bht_value; // @[Frontend.scala 273:35 Frontend.scala 273:35]
  assign btb_io_ras_update_valid = taken_idx ? _T_598 : _T_331; // @[Frontend.scala 187:29 Frontend.scala 250:33 Frontend.scala 250:33]
  assign btb_io_ras_update_bits_cfiType = taken_idx ? _T_606 : _T_339; // @[Frontend.scala 251:40 Frontend.scala 251:40]
  assign btb_io_ras_update_bits_returnAddr = _T_103[38:0]; // @[Frontend.scala 304:39]
  assign btb_io_flush = _T_588 | _T_321; // @[Frontend.scala 182:18 Frontend.scala 200:54 Frontend.scala 241:22 Frontend.scala 241:22]
  assign Frontend_cov_read_addr = Frontend_state;
  assign Frontend_cov_read_data = Frontend_cov[Frontend_cov_read_addr]; // @[Coverage map for Frontend]
  assign Frontend_cov_write_data = 1'h1;
  assign Frontend_cov_write_addr = Frontend_state;
  assign Frontend_cov_write_mask = 1'h1;
  assign Frontend_cov_write_en = 1'h1;
  assign s2_partial_insn_valid_shl = s2_partial_insn_valid;
  assign s2_partial_insn_valid_pad = {5'h0,s2_partial_insn_valid_shl};
  assign _T_37_shl = {_T_37, 1'h0};
  assign _T_37_pad = {4'h0,_T_37_shl};
  assign s2_btb_resp_valid_shl = {s2_btb_resp_valid, 2'h0};
  assign s2_btb_resp_valid_pad = {3'h0,s2_btb_resp_valid_shl};
  assign s2_btb_resp_bits_taken_shl = {s2_btb_resp_bits_taken, 3'h0};
  assign s2_btb_resp_bits_taken_pad = {2'h0,s2_btb_resp_bits_taken_shl};
  assign s2_btb_resp_bits_bht_value_shl = {s2_btb_resp_bits_bht_value, 4'h0};
  assign s2_btb_resp_bits_bht_value_pad = {1'h0,s2_btb_resp_bits_bht_value_shl};
  assign s2_valid_shl = {s2_valid, 5'h0};
  assign s2_valid_pad = s2_valid_shl;
  assign Frontend_xor4 = _T_37_pad ^ s2_btb_resp_valid_pad;
  assign Frontend_xor1 = s2_partial_insn_valid_pad ^ Frontend_xor4;
  assign Frontend_xor6 = s2_btb_resp_bits_bht_value_pad ^ s2_valid_pad;
  assign Frontend_xor2 = s2_btb_resp_bits_taken_pad ^ Frontend_xor6;
  assign Frontend_xor0 = Frontend_xor1 ^ Frontend_xor2;
  assign icache_sum = Frontend_covSum + icache_io_covSum;
  assign fq_sum = icache_sum + fq_io_covSum;
  assign tlb_sum = fq_sum + tlb_io_covSum;
  assign btb_sum = tlb_sum + btb_io_covSum;
  assign io_covSum = btb_sum;
  assign stopEn0 = ~_T_9;
  assign stopEn1 = ~_T_82;
  assign stopEn2 = ~_T_654;
  assign icache_metaAssert_wire = icache_metaAssert;
  assign fq_metaAssert_wire = fq_metaAssert;
  assign tlb_metaAssert_wire = tlb_metaAssert;
  assign btb_metaAssert_wire = btb_metaAssert;
  assign Frontend_or4 = stopEn1 | stopEn2;
  assign Frontend_or1 = stopEn0 | Frontend_or4;
  assign Frontend_or5 = icache_metaAssert_wire | fq_metaAssert_wire;
  assign Frontend_or6 = tlb_metaAssert_wire | btb_metaAssert_wire;
  assign Frontend_or2 = Frontend_or5 | Frontend_or6;
  assign Frontend_or0 = Frontend_or1 | Frontend_or2;
  assign metaAssert = Frontend_or0;
  assign icache_metaReset = metaReset | icache_halt;
  assign fq_metaReset = metaReset | fq_halt;
  assign tlb_metaReset = metaReset | tlb_halt;
  assign btb_metaReset = metaReset | btb_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  s2_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  s1_pc = _RAND_2[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  s1_speculative = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  s2_pc = _RAND_4[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  s2_btb_resp_valid = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  s2_btb_resp_bits_taken = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  s2_btb_resp_bits_bridx = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  s2_btb_resp_bits_entry = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  s2_btb_resp_bits_bht_history = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  s2_btb_resp_bits_bht_value = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  s2_tlb_resp_miss = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  s2_tlb_resp_pf_inst = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  s2_tlb_resp_ae_inst = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  s2_tlb_resp_cacheable = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  s2_speculative = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  s2_partial_insn_valid = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  s2_partial_insn = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  wrong_path = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_37 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_59 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  Frontend_state = _RAND_21[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    Frontend_cov[initvar] = _RAND_22[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  Frontend_covSum = _RAND_23[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge gated_clock) begin
    if (metaReset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= io_cpu_req_valid | s0_fq_has_space;
    end
    if (metaReset) begin
      s2_valid <= 1'h0;
    end else if (reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= _GEN_0;
    end
    if (metaReset) begin
      s1_pc <= 40'h0;
    end else begin
      s1_pc <= io_cpu_npc;
    end
    if (metaReset) begin
      s1_speculative <= 1'h0;
    end else if (io_cpu_req_valid) begin
      s1_speculative <= io_cpu_req_bits_speculative;
    end else if (s2_replay) begin
      s1_speculative <= s2_speculative;
    end else begin
      s1_speculative <= s0_speculative;
    end
    if (metaReset) begin
      s2_pc <= 40'h0;
    end else if (reset) begin
      s2_pc <= {{8'd0}, ~_T_27};
    end else if (~s2_replay) begin
      s2_pc <= s1_pc;
    end
    if (metaReset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if (metaReset) begin
      s2_btb_resp_bits_taken <= 1'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if (metaReset) begin
      s2_btb_resp_bits_bridx <= 1'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_bridx <= btb_io_resp_bits_bridx;
    end
    if (metaReset) begin
      s2_btb_resp_bits_entry <= 5'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if (metaReset) begin
      s2_btb_resp_bits_bht_history <= 8'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_bht_history <= btb_io_resp_bits_bht_history;
    end
    if (metaReset) begin
      s2_btb_resp_bits_bht_value <= 1'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if (metaReset) begin
      s2_tlb_resp_miss <= 1'h0;
    end else if (~s2_replay) begin
      s2_tlb_resp_miss <= tlb_io_resp_miss;
    end
    if (metaReset) begin
      s2_tlb_resp_pf_inst <= 1'h0;
    end else if (~s2_replay) begin
      s2_tlb_resp_pf_inst <= tlb_io_resp_pf_inst;
    end
    if (metaReset) begin
      s2_tlb_resp_ae_inst <= 1'h0;
    end else if (~s2_replay) begin
      s2_tlb_resp_ae_inst <= tlb_io_resp_ae_inst;
    end
    if (metaReset) begin
      s2_tlb_resp_cacheable <= 1'h0;
    end else if (~s2_replay) begin
      s2_tlb_resp_cacheable <= tlb_io_resp_cacheable;
    end
    if (metaReset) begin
      s2_speculative <= 1'h0;
    end else if (reset) begin
      s2_speculative <= 1'h0;
    end else if (~s2_replay) begin
      s2_speculative <= s1_speculative;
    end
    if (metaReset) begin
      s2_partial_insn_valid <= 1'h0;
    end else if (reset) begin
      s2_partial_insn_valid <= 1'h0;
    end else if (s2_redirect) begin
      s2_partial_insn_valid <= 1'h0;
    end else if (_T_647) begin
      s2_partial_insn_valid <= 1'h0;
    end else if (_T_32) begin
      s2_partial_insn_valid <= _T_643;
    end
    if (metaReset) begin
      s2_partial_insn <= 16'h0;
    end else if (_T_32) begin
      if (_T_643) begin
        s2_partial_insn <= _T_644;
      end
    end
    if (metaReset) begin
      wrong_path <= 1'h0;
    end else if (io_cpu_req_valid) begin
      wrong_path <= 1'h0;
    end else if (taken_idx) begin
      if (~s2_btb_taken) begin
        wrong_path <= _GEN_77;
      end else begin
        wrong_path <= _GEN_76;
      end
    end else begin
      wrong_path <= _GEN_76;
    end
    if (metaReset) begin
      _T_37 <= 1'h0;
    end else begin
      _T_37 <= reset | _T_36;
    end
    if (metaReset) begin
      _T_59 <= 1'h0;
    end else begin
      _T_59 <= s1_valid;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_9) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Frontend.scala:91 assert(!(io.cpu.req.valid || io.cpu.sfence.valid || io.cpu.flush_icache || io.cpu.bht_update.valid || io.cpu.btb_update.valid) || io.cpu.might_request)\n"); // @[Frontend.scala 91:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_9) begin
          $fatal; // @[Frontend.scala 91:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_82) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Frontend.scala:177 assert(!(s2_speculative && io.ptw.customCSRs.asInstanceOf[RocketCustomCSRs].disableSpeculativeICacheRefill && !icache.io.s2_kill))\n"); // @[Frontend.scala 177:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_82) begin
          $fatal; // @[Frontend.scala 177:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_654) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Frontend.scala:322 assert(!s2_partial_insn_valid || fq.io.enq.bits.mask(0))\n"); // @[Frontend.scala 322:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_654) begin
          $fatal; // @[Frontend.scala 322:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    Frontend_state <= Frontend_xor0;
    if (!(Frontend_cov_read_data)) begin
      Frontend_covSum <= Frontend_covSum + 1'h1;
    end
  end
  always @(posedge gated_clock) begin
    if(Frontend_cov_write_en & Frontend_cov_write_mask) begin
      Frontend_cov[Frontend_cov_write_addr] <= Frontend_cov_write_data; // @[Coverage map for Frontend]
    end
  end
endmodule
module TLBuffer_7(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [3:0]  auto_in_a_bits_size,
  input  [1:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_a_bits_corrupt,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [2:0]  auto_in_b_bits_opcode,
  output [1:0]  auto_in_b_bits_param,
  output [3:0]  auto_in_b_bits_size,
  output [1:0]  auto_in_b_bits_source,
  output [31:0] auto_in_b_bits_address,
  output [7:0]  auto_in_b_bits_mask,
  output        auto_in_b_bits_corrupt,
  output        auto_in_c_ready,
  input         auto_in_c_valid,
  input  [2:0]  auto_in_c_bits_opcode,
  input  [2:0]  auto_in_c_bits_param,
  input  [3:0]  auto_in_c_bits_size,
  input  [1:0]  auto_in_c_bits_source,
  input  [31:0] auto_in_c_bits_address,
  input  [63:0] auto_in_c_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [3:0]  auto_in_d_bits_size,
  output [1:0]  auto_in_d_bits_source,
  output [1:0]  auto_in_d_bits_sink,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  output        auto_in_e_ready,
  input         auto_in_e_valid,
  input  [1:0]  auto_in_e_bits_sink,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [1:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_a_bits_corrupt,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [2:0]  auto_out_b_bits_opcode,
  input  [1:0]  auto_out_b_bits_param,
  input  [3:0]  auto_out_b_bits_size,
  input  [1:0]  auto_out_b_bits_source,
  input  [31:0] auto_out_b_bits_address,
  input  [7:0]  auto_out_b_bits_mask,
  input         auto_out_b_bits_corrupt,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [3:0]  auto_out_c_bits_size,
  output [1:0]  auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output        auto_out_c_bits_corrupt,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [3:0]  auto_out_d_bits_size,
  input  [1:0]  auto_out_d_bits_source,
  input  [1:0]  auto_out_d_bits_sink,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output [1:0]  auto_out_e_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         Queue_3_halt,
  input         Queue_halt,
  input         TLMonitor_halt,
  input         Queue_2_halt,
  input         Queue_4_halt,
  input         Queue_1_halt
);
  wire  TLMonitor_clock; // @[Nodes.scala 25:25]
  wire  TLMonitor_reset; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_a_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_a_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_a_bits_opcode; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_a_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_a_bits_size; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_a_bits_source; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_io_in_a_bits_address; // @[Nodes.scala 25:25]
  wire [7:0] TLMonitor_io_in_a_bits_mask; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_a_bits_corrupt; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_b_bits_opcode; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_b_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_b_bits_size; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_b_bits_source; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_io_in_b_bits_address; // @[Nodes.scala 25:25]
  wire [7:0] TLMonitor_io_in_b_bits_mask; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_bits_corrupt; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_c_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_c_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_c_bits_opcode; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_c_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_c_bits_size; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_c_bits_source; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_io_in_c_bits_address; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_d_bits_opcode; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_d_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_d_bits_size; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_d_bits_source; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_d_bits_sink; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_bits_denied; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_bits_corrupt; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_e_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_e_valid; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_e_bits_sink; // @[Nodes.scala 25:25]
  wire [29:0] TLMonitor_io_covSum; // @[Nodes.scala 25:25]
  wire  TLMonitor_metaAssert; // @[Nodes.scala 25:25]
  wire  TLMonitor_metaReset; // @[Nodes.scala 25:25]
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_io_enq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_io_enq_bits_param; // @[Decoupled.scala 296:21]
  wire [3:0] Queue_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_io_enq_bits_source; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_address; // @[Decoupled.scala 296:21]
  wire [7:0] Queue_io_enq_bits_mask; // @[Decoupled.scala 296:21]
  wire [63:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_corrupt; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_io_deq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_io_deq_bits_param; // @[Decoupled.scala 296:21]
  wire [3:0] Queue_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_io_deq_bits_source; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_address; // @[Decoupled.scala 296:21]
  wire [7:0] Queue_io_deq_bits_mask; // @[Decoupled.scala 296:21]
  wire [63:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_corrupt; // @[Decoupled.scala 296:21]
  wire [29:0] Queue_io_covSum; // @[Decoupled.scala 296:21]
  wire  Queue_metaAssert; // @[Decoupled.scala 296:21]
  wire  Queue_metaReset; // @[Decoupled.scala 296:21]
  wire  Queue_1_clock; // @[Decoupled.scala 296:21]
  wire  Queue_1_reset; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_1_io_enq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_1_io_enq_bits_param; // @[Decoupled.scala 296:21]
  wire [3:0] Queue_1_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_1_io_enq_bits_source; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_1_io_enq_bits_sink; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_enq_bits_denied; // @[Decoupled.scala 296:21]
  wire [63:0] Queue_1_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_enq_bits_corrupt; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_1_io_deq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_1_io_deq_bits_param; // @[Decoupled.scala 296:21]
  wire [3:0] Queue_1_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_1_io_deq_bits_source; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_1_io_deq_bits_sink; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_deq_bits_denied; // @[Decoupled.scala 296:21]
  wire [63:0] Queue_1_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_deq_bits_corrupt; // @[Decoupled.scala 296:21]
  wire [29:0] Queue_1_io_covSum; // @[Decoupled.scala 296:21]
  wire  Queue_1_metaAssert; // @[Decoupled.scala 296:21]
  wire  Queue_1_metaReset; // @[Decoupled.scala 296:21]
  wire  Queue_2_clock; // @[Decoupled.scala 296:21]
  wire  Queue_2_reset; // @[Decoupled.scala 296:21]
  wire  Queue_2_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_2_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_2_io_enq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_2_io_enq_bits_param; // @[Decoupled.scala 296:21]
  wire [3:0] Queue_2_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_2_io_enq_bits_source; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_2_io_enq_bits_address; // @[Decoupled.scala 296:21]
  wire [7:0] Queue_2_io_enq_bits_mask; // @[Decoupled.scala 296:21]
  wire  Queue_2_io_enq_bits_corrupt; // @[Decoupled.scala 296:21]
  wire  Queue_2_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_2_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_2_io_deq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_2_io_deq_bits_param; // @[Decoupled.scala 296:21]
  wire [3:0] Queue_2_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_2_io_deq_bits_source; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_2_io_deq_bits_address; // @[Decoupled.scala 296:21]
  wire [7:0] Queue_2_io_deq_bits_mask; // @[Decoupled.scala 296:21]
  wire  Queue_2_io_deq_bits_corrupt; // @[Decoupled.scala 296:21]
  wire [29:0] Queue_2_io_covSum; // @[Decoupled.scala 296:21]
  wire  Queue_2_metaAssert; // @[Decoupled.scala 296:21]
  wire  Queue_2_metaReset; // @[Decoupled.scala 296:21]
  wire  Queue_3_clock; // @[Decoupled.scala 296:21]
  wire  Queue_3_reset; // @[Decoupled.scala 296:21]
  wire  Queue_3_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_3_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_3_io_enq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_3_io_enq_bits_param; // @[Decoupled.scala 296:21]
  wire [3:0] Queue_3_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_3_io_enq_bits_source; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_3_io_enq_bits_address; // @[Decoupled.scala 296:21]
  wire [63:0] Queue_3_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_3_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_3_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_3_io_deq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_3_io_deq_bits_param; // @[Decoupled.scala 296:21]
  wire [3:0] Queue_3_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_3_io_deq_bits_source; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_3_io_deq_bits_address; // @[Decoupled.scala 296:21]
  wire [63:0] Queue_3_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_3_io_deq_bits_corrupt; // @[Decoupled.scala 296:21]
  wire [29:0] Queue_3_io_covSum; // @[Decoupled.scala 296:21]
  wire  Queue_3_metaAssert; // @[Decoupled.scala 296:21]
  wire  Queue_3_metaReset; // @[Decoupled.scala 296:21]
  wire  Queue_4_clock; // @[Decoupled.scala 296:21]
  wire  Queue_4_reset; // @[Decoupled.scala 296:21]
  wire  Queue_4_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_4_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_4_io_enq_bits_sink; // @[Decoupled.scala 296:21]
  wire  Queue_4_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_4_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_4_io_deq_bits_sink; // @[Decoupled.scala 296:21]
  wire [29:0] Queue_4_io_covSum; // @[Decoupled.scala 296:21]
  wire  Queue_4_metaAssert; // @[Decoupled.scala 296:21]
  wire  Queue_4_metaReset; // @[Decoupled.scala 296:21]
  wire [29:0] TLBuffer_7_covSum;
  wire [29:0] Queue_3_sum;
  wire [29:0] Queue_sum;
  wire [29:0] TLMonitor_sum;
  wire [29:0] Queue_2_sum;
  wire [29:0] Queue_4_sum;
  wire [29:0] Queue_1_sum;
  wire  TLMonitor_metaAssert_wire;
  wire  Queue_metaAssert_wire;
  wire  Queue_1_metaAssert_wire;
  wire  Queue_4_metaAssert_wire;
  wire  Queue_3_metaAssert_wire;
  wire  Queue_2_metaAssert_wire;
  wire  TLBuffer_7_or4;
  wire  TLBuffer_7_or1;
  wire  TLBuffer_7_or6;
  wire  TLBuffer_7_or2;
  wire  TLBuffer_7_or0;
  reg  TLBuffer_7_metaAssert;
  reg [31:0] _RAND_0;
  TLMonitor_37 TLMonitor ( // @[Nodes.scala 25:25]
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_b_ready(TLMonitor_io_in_b_ready),
    .io_in_b_valid(TLMonitor_io_in_b_valid),
    .io_in_b_bits_opcode(TLMonitor_io_in_b_bits_opcode),
    .io_in_b_bits_param(TLMonitor_io_in_b_bits_param),
    .io_in_b_bits_size(TLMonitor_io_in_b_bits_size),
    .io_in_b_bits_source(TLMonitor_io_in_b_bits_source),
    .io_in_b_bits_address(TLMonitor_io_in_b_bits_address),
    .io_in_b_bits_mask(TLMonitor_io_in_b_bits_mask),
    .io_in_b_bits_corrupt(TLMonitor_io_in_b_bits_corrupt),
    .io_in_c_ready(TLMonitor_io_in_c_ready),
    .io_in_c_valid(TLMonitor_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_io_in_c_bits_address),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt),
    .io_in_e_ready(TLMonitor_io_in_e_ready),
    .io_in_e_valid(TLMonitor_io_in_e_valid),
    .io_in_e_bits_sink(TLMonitor_io_in_e_bits_sink),
    .io_covSum(TLMonitor_io_covSum),
    .metaAssert(TLMonitor_metaAssert),
    .metaReset(TLMonitor_metaReset)
  );
  Queue_32 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_opcode(Queue_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_io_enq_bits_param),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_source(Queue_io_enq_bits_source),
    .io_enq_bits_address(Queue_io_enq_bits_address),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_corrupt(Queue_io_enq_bits_corrupt),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_io_deq_bits_param),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source),
    .io_deq_bits_address(Queue_io_deq_bits_address),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_corrupt(Queue_io_deq_bits_corrupt),
    .io_covSum(Queue_io_covSum),
    .metaAssert(Queue_metaAssert),
    .metaReset(Queue_metaReset)
  );
  Queue_33 Queue_1 ( // @[Decoupled.scala 296:21]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_opcode(Queue_1_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_1_io_enq_bits_param),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_source(Queue_1_io_enq_bits_source),
    .io_enq_bits_sink(Queue_1_io_enq_bits_sink),
    .io_enq_bits_denied(Queue_1_io_enq_bits_denied),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_corrupt(Queue_1_io_enq_bits_corrupt),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_opcode(Queue_1_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_1_io_deq_bits_param),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_source(Queue_1_io_deq_bits_source),
    .io_deq_bits_sink(Queue_1_io_deq_bits_sink),
    .io_deq_bits_denied(Queue_1_io_deq_bits_denied),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_corrupt(Queue_1_io_deq_bits_corrupt),
    .io_covSum(Queue_1_io_covSum),
    .metaAssert(Queue_1_metaAssert),
    .metaReset(Queue_1_metaReset)
  );
  Queue_34 Queue_2 ( // @[Decoupled.scala 296:21]
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_opcode(Queue_2_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_2_io_enq_bits_param),
    .io_enq_bits_size(Queue_2_io_enq_bits_size),
    .io_enq_bits_source(Queue_2_io_enq_bits_source),
    .io_enq_bits_address(Queue_2_io_enq_bits_address),
    .io_enq_bits_mask(Queue_2_io_enq_bits_mask),
    .io_enq_bits_corrupt(Queue_2_io_enq_bits_corrupt),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_opcode(Queue_2_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_2_io_deq_bits_param),
    .io_deq_bits_size(Queue_2_io_deq_bits_size),
    .io_deq_bits_source(Queue_2_io_deq_bits_source),
    .io_deq_bits_address(Queue_2_io_deq_bits_address),
    .io_deq_bits_mask(Queue_2_io_deq_bits_mask),
    .io_deq_bits_corrupt(Queue_2_io_deq_bits_corrupt),
    .io_covSum(Queue_2_io_covSum),
    .metaAssert(Queue_2_metaAssert),
    .metaReset(Queue_2_metaReset)
  );
  Queue_35 Queue_3 ( // @[Decoupled.scala 296:21]
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_opcode(Queue_3_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_3_io_enq_bits_param),
    .io_enq_bits_size(Queue_3_io_enq_bits_size),
    .io_enq_bits_source(Queue_3_io_enq_bits_source),
    .io_enq_bits_address(Queue_3_io_enq_bits_address),
    .io_enq_bits_data(Queue_3_io_enq_bits_data),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_opcode(Queue_3_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_3_io_deq_bits_param),
    .io_deq_bits_size(Queue_3_io_deq_bits_size),
    .io_deq_bits_source(Queue_3_io_deq_bits_source),
    .io_deq_bits_address(Queue_3_io_deq_bits_address),
    .io_deq_bits_data(Queue_3_io_deq_bits_data),
    .io_deq_bits_corrupt(Queue_3_io_deq_bits_corrupt),
    .io_covSum(Queue_3_io_covSum),
    .metaAssert(Queue_3_metaAssert),
    .metaReset(Queue_3_metaReset)
  );
  Queue_36 Queue_4 ( // @[Decoupled.scala 296:21]
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_sink(Queue_4_io_enq_bits_sink),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_sink(Queue_4_io_deq_bits_sink),
    .io_covSum(Queue_4_io_covSum),
    .metaAssert(Queue_4_metaAssert),
    .metaReset(Queue_4_metaReset)
  );
  assign auto_in_a_ready = Queue_io_enq_ready; // @[LazyModule.scala 303:16]
  assign auto_in_b_valid = Queue_2_io_deq_valid; // @[LazyModule.scala 303:16]
  assign auto_in_b_bits_opcode = Queue_2_io_deq_bits_opcode; // @[LazyModule.scala 303:16]
  assign auto_in_b_bits_param = Queue_2_io_deq_bits_param; // @[LazyModule.scala 303:16]
  assign auto_in_b_bits_size = Queue_2_io_deq_bits_size; // @[LazyModule.scala 303:16]
  assign auto_in_b_bits_source = Queue_2_io_deq_bits_source; // @[LazyModule.scala 303:16]
  assign auto_in_b_bits_address = Queue_2_io_deq_bits_address; // @[LazyModule.scala 303:16]
  assign auto_in_b_bits_mask = Queue_2_io_deq_bits_mask; // @[LazyModule.scala 303:16]
  assign auto_in_b_bits_corrupt = Queue_2_io_deq_bits_corrupt; // @[LazyModule.scala 303:16]
  assign auto_in_c_ready = Queue_3_io_enq_ready; // @[LazyModule.scala 303:16]
  assign auto_in_d_valid = Queue_1_io_deq_valid; // @[LazyModule.scala 303:16]
  assign auto_in_d_bits_opcode = Queue_1_io_deq_bits_opcode; // @[LazyModule.scala 303:16]
  assign auto_in_d_bits_param = Queue_1_io_deq_bits_param; // @[LazyModule.scala 303:16]
  assign auto_in_d_bits_size = Queue_1_io_deq_bits_size; // @[LazyModule.scala 303:16]
  assign auto_in_d_bits_source = Queue_1_io_deq_bits_source; // @[LazyModule.scala 303:16]
  assign auto_in_d_bits_sink = Queue_1_io_deq_bits_sink; // @[LazyModule.scala 303:16]
  assign auto_in_d_bits_denied = Queue_1_io_deq_bits_denied; // @[LazyModule.scala 303:16]
  assign auto_in_d_bits_data = Queue_1_io_deq_bits_data; // @[LazyModule.scala 303:16]
  assign auto_in_d_bits_corrupt = Queue_1_io_deq_bits_corrupt; // @[LazyModule.scala 303:16]
  assign auto_in_e_ready = Queue_4_io_enq_ready; // @[LazyModule.scala 303:16]
  assign auto_out_a_valid = Queue_io_deq_valid; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_opcode = Queue_io_deq_bits_opcode; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_param = Queue_io_deq_bits_param; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_size = Queue_io_deq_bits_size; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_source = Queue_io_deq_bits_source; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_address = Queue_io_deq_bits_address; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_mask = Queue_io_deq_bits_mask; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 305:12]
  assign auto_out_a_bits_corrupt = Queue_io_deq_bits_corrupt; // @[LazyModule.scala 305:12]
  assign auto_out_b_ready = Queue_2_io_enq_ready; // @[LazyModule.scala 305:12]
  assign auto_out_c_valid = Queue_3_io_deq_valid; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_opcode = Queue_3_io_deq_bits_opcode; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_param = Queue_3_io_deq_bits_param; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_size = Queue_3_io_deq_bits_size; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_source = Queue_3_io_deq_bits_source; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_address = Queue_3_io_deq_bits_address; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_data = Queue_3_io_deq_bits_data; // @[LazyModule.scala 305:12]
  assign auto_out_c_bits_corrupt = Queue_3_io_deq_bits_corrupt; // @[LazyModule.scala 305:12]
  assign auto_out_d_ready = Queue_1_io_enq_ready; // @[LazyModule.scala 305:12]
  assign auto_out_e_valid = Queue_4_io_deq_valid; // @[LazyModule.scala 305:12]
  assign auto_out_e_bits_sink = Queue_4_io_deq_bits_sink; // @[LazyModule.scala 305:12]
  assign TLMonitor_clock = clock;
  assign TLMonitor_reset = reset;
  assign TLMonitor_io_in_a_ready = Queue_io_enq_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_ready = auto_in_b_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_valid = Queue_2_io_deq_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_opcode = Queue_2_io_deq_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_param = Queue_2_io_deq_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_size = Queue_2_io_deq_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_source = Queue_2_io_deq_bits_source; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_address = Queue_2_io_deq_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_mask = Queue_2_io_deq_bits_mask; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_corrupt = Queue_2_io_deq_bits_corrupt; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_ready = Queue_3_io_enq_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_valid = auto_in_c_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_source = auto_in_c_bits_source; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_valid = Queue_1_io_deq_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_opcode = Queue_1_io_deq_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_param = Queue_1_io_deq_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_size = Queue_1_io_deq_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_source = Queue_1_io_deq_bits_source; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_sink = Queue_1_io_deq_bits_sink; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_denied = Queue_1_io_deq_bits_denied; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_corrupt = Queue_1_io_deq_bits_corrupt; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_e_ready = Queue_4_io_enq_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_e_valid = auto_in_e_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_e_bits_sink = auto_in_e_bits_sink; // @[Nodes.scala 26:19]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_a_valid; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_param = auto_in_a_bits_param; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_size = auto_in_a_bits_size; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_source = auto_in_a_bits_source; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_address = auto_in_a_bits_address; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_mask = auto_in_a_bits_mask; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = auto_in_a_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = auto_out_a_ready; // @[Buffer.scala 38:13]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = auto_out_d_valid; // @[Decoupled.scala 297:22]
  assign Queue_1_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Decoupled.scala 298:21]
  assign Queue_1_io_enq_bits_param = auto_out_d_bits_param; // @[Decoupled.scala 298:21]
  assign Queue_1_io_enq_bits_size = auto_out_d_bits_size; // @[Decoupled.scala 298:21]
  assign Queue_1_io_enq_bits_source = auto_out_d_bits_source; // @[Decoupled.scala 298:21]
  assign Queue_1_io_enq_bits_sink = auto_out_d_bits_sink; // @[Decoupled.scala 298:21]
  assign Queue_1_io_enq_bits_denied = auto_out_d_bits_denied; // @[Decoupled.scala 298:21]
  assign Queue_1_io_enq_bits_data = auto_out_d_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_1_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Decoupled.scala 298:21]
  assign Queue_1_io_deq_ready = auto_in_d_ready; // @[Buffer.scala 39:13]
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = auto_out_b_valid; // @[Decoupled.scala 297:22]
  assign Queue_2_io_enq_bits_opcode = auto_out_b_bits_opcode; // @[Decoupled.scala 298:21]
  assign Queue_2_io_enq_bits_param = auto_out_b_bits_param; // @[Decoupled.scala 298:21]
  assign Queue_2_io_enq_bits_size = auto_out_b_bits_size; // @[Decoupled.scala 298:21]
  assign Queue_2_io_enq_bits_source = auto_out_b_bits_source; // @[Decoupled.scala 298:21]
  assign Queue_2_io_enq_bits_address = auto_out_b_bits_address; // @[Decoupled.scala 298:21]
  assign Queue_2_io_enq_bits_mask = auto_out_b_bits_mask; // @[Decoupled.scala 298:21]
  assign Queue_2_io_enq_bits_corrupt = auto_out_b_bits_corrupt; // @[Decoupled.scala 298:21]
  assign Queue_2_io_deq_ready = auto_in_b_ready; // @[Buffer.scala 42:15]
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = auto_in_c_valid; // @[Decoupled.scala 297:22]
  assign Queue_3_io_enq_bits_opcode = auto_in_c_bits_opcode; // @[Decoupled.scala 298:21]
  assign Queue_3_io_enq_bits_param = auto_in_c_bits_param; // @[Decoupled.scala 298:21]
  assign Queue_3_io_enq_bits_size = auto_in_c_bits_size; // @[Decoupled.scala 298:21]
  assign Queue_3_io_enq_bits_source = auto_in_c_bits_source; // @[Decoupled.scala 298:21]
  assign Queue_3_io_enq_bits_address = auto_in_c_bits_address; // @[Decoupled.scala 298:21]
  assign Queue_3_io_enq_bits_data = auto_in_c_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_3_io_deq_ready = auto_out_c_ready; // @[Buffer.scala 43:15]
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = auto_in_e_valid; // @[Decoupled.scala 297:22]
  assign Queue_4_io_enq_bits_sink = auto_in_e_bits_sink; // @[Decoupled.scala 298:21]
  assign Queue_4_io_deq_ready = auto_out_e_ready; // @[Buffer.scala 44:15]
  assign TLBuffer_7_covSum = 30'h0;
  assign Queue_3_sum = TLBuffer_7_covSum + Queue_3_io_covSum;
  assign Queue_sum = Queue_3_sum + Queue_io_covSum;
  assign TLMonitor_sum = Queue_sum + TLMonitor_io_covSum;
  assign Queue_2_sum = TLMonitor_sum + Queue_2_io_covSum;
  assign Queue_4_sum = Queue_2_sum + Queue_4_io_covSum;
  assign Queue_1_sum = Queue_4_sum + Queue_1_io_covSum;
  assign io_covSum = Queue_1_sum;
  assign TLMonitor_metaAssert_wire = TLMonitor_metaAssert;
  assign Queue_2_metaAssert_wire = Queue_2_metaAssert;
  assign Queue_4_metaAssert_wire = Queue_4_metaAssert;
  assign Queue_1_metaAssert_wire = Queue_1_metaAssert;
  assign Queue_metaAssert_wire = Queue_metaAssert;
  assign Queue_3_metaAssert_wire = Queue_3_metaAssert;
  assign TLBuffer_7_or4 = Queue_4_metaAssert_wire | TLMonitor_metaAssert_wire;
  assign TLBuffer_7_or1 = Queue_2_metaAssert_wire | TLBuffer_7_or4;
  assign TLBuffer_7_or6 = Queue_metaAssert_wire | Queue_3_metaAssert_wire;
  assign TLBuffer_7_or2 = Queue_1_metaAssert_wire | TLBuffer_7_or6;
  assign TLBuffer_7_or0 = TLBuffer_7_or1 | TLBuffer_7_or2;
  assign metaAssert = TLBuffer_7_metaAssert;
  assign Queue_3_metaReset = metaReset | Queue_3_halt;
  assign Queue_metaReset = metaReset | Queue_halt;
  assign TLMonitor_metaReset = metaReset | TLMonitor_halt;
  assign Queue_2_metaReset = metaReset | Queue_2_halt;
  assign Queue_4_metaReset = metaReset | Queue_4_halt;
  assign Queue_1_metaReset = metaReset | Queue_1_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  TLBuffer_7_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      TLBuffer_7_metaAssert <= 1'h0;
    end else begin
      TLBuffer_7_metaAssert <= TLBuffer_7_metaAssert | TLBuffer_7_or0;
    end
  end
endmodule
module IntSyncAsyncCrossingSink(
  input         clock,
  input         auto_in_sync_0,
  output        auto_out_0,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         SynchronizerShiftReg_w1_d3_halt
);
  wire  SynchronizerShiftReg_w1_d3_clock; // @[ShiftReg.scala 45:23]
  wire  SynchronizerShiftReg_w1_d3_io_d; // @[ShiftReg.scala 45:23]
  wire  SynchronizerShiftReg_w1_d3_io_q; // @[ShiftReg.scala 45:23]
  wire [29:0] SynchronizerShiftReg_w1_d3_io_covSum; // @[ShiftReg.scala 45:23]
  wire  SynchronizerShiftReg_w1_d3_metaAssert; // @[ShiftReg.scala 45:23]
  wire  SynchronizerShiftReg_w1_d3_metaReset; // @[ShiftReg.scala 45:23]
  wire  SynchronizerShiftReg_w1_d3_NonSyncResetSynchronizerPrimitiveShiftReg_d3_halt; // @[ShiftReg.scala 45:23]
  wire [29:0] IntSyncAsyncCrossingSink_covSum;
  wire [29:0] SynchronizerShiftReg_w1_d3_sum;
  wire  SynchronizerShiftReg_w1_d3_metaAssert_wire;
  SynchronizerShiftReg_w1_d3 SynchronizerShiftReg_w1_d3 ( // @[ShiftReg.scala 45:23]
    .clock(SynchronizerShiftReg_w1_d3_clock),
    .io_d(SynchronizerShiftReg_w1_d3_io_d),
    .io_q(SynchronizerShiftReg_w1_d3_io_q),
    .io_covSum(SynchronizerShiftReg_w1_d3_io_covSum),
    .metaAssert(SynchronizerShiftReg_w1_d3_metaAssert),
    .metaReset(SynchronizerShiftReg_w1_d3_metaReset),
    .NonSyncResetSynchronizerPrimitiveShiftReg_d3_halt(SynchronizerShiftReg_w1_d3_NonSyncResetSynchronizerPrimitiveShiftReg_d3_halt)
  );
  assign auto_out_0 = SynchronizerShiftReg_w1_d3_io_q; // @[LazyModule.scala 305:12]
  assign SynchronizerShiftReg_w1_d3_clock = clock;
  assign SynchronizerShiftReg_w1_d3_io_d = auto_in_sync_0; // @[ShiftReg.scala 47:16]
  assign IntSyncAsyncCrossingSink_covSum = 30'h0;
  assign SynchronizerShiftReg_w1_d3_sum = IntSyncAsyncCrossingSink_covSum + SynchronizerShiftReg_w1_d3_io_covSum;
  assign io_covSum = SynchronizerShiftReg_w1_d3_sum;
  assign SynchronizerShiftReg_w1_d3_metaAssert_wire = SynchronizerShiftReg_w1_d3_metaAssert;
  assign metaAssert = SynchronizerShiftReg_w1_d3_metaAssert_wire;
  assign SynchronizerShiftReg_w1_d3_metaReset = metaReset | SynchronizerShiftReg_w1_d3_halt;
endmodule
module IntSyncSyncCrossingSink(
  input         auto_in_sync_0,
  input         auto_in_sync_1,
  output        auto_out_0,
  output        auto_out_1,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] IntSyncSyncCrossingSink_covSum;
  assign auto_out_0 = auto_in_sync_0; // @[LazyModule.scala 305:12]
  assign auto_out_1 = auto_in_sync_1; // @[LazyModule.scala 305:12]
  assign IntSyncSyncCrossingSink_covSum = 30'h0;
  assign io_covSum = IntSyncSyncCrossingSink_covSum;
  assign metaAssert = 1'h0;
endmodule
module IntSyncSyncCrossingSink_1(
  input         auto_in_sync_0,
  output        auto_out_0,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] IntSyncSyncCrossingSink_1_covSum;
  assign auto_out_0 = auto_in_sync_0; // @[LazyModule.scala 305:12]
  assign IntSyncSyncCrossingSink_1_covSum = 30'h0;
  assign io_covSum = IntSyncSyncCrossingSink_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module FPU(
  input         clock,
  input         reset,
  input  [31:0] io_inst,
  input  [63:0] io_fromint_data,
  input  [2:0]  io_fcsr_rm,
  output        io_fcsr_flags_valid,
  output [4:0]  io_fcsr_flags_bits,
  output [63:0] io_store_data,
  output [63:0] io_toint_data,
  input         io_dmem_resp_val,
  input  [2:0]  io_dmem_resp_type,
  input  [4:0]  io_dmem_resp_tag,
  input  [63:0] io_dmem_resp_data,
  input         io_valid,
  output        io_fcsr_rdy,
  output        io_nack_mem,
  output        io_illegal_rm,
  input         io_killx,
  input         io_killm,
  output        io_dec_wen,
  output        io_dec_ren1,
  output        io_dec_ren2,
  output        io_dec_ren3,
  output        io_sboard_set,
  output        io_sboard_clr,
  output [4:0]  io_sboard_clra,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         divSqrt_1_halt,
  input         ifpu_halt,
  input         divSqrt_halt,
  input         fpmu_halt,
  input         dfma_halt,
  input         fpiu_halt,
  input         sfma_halt,
  output [19:0] Checking_FPU_regstate,	//Jaewon_FPU_regstate
  output [29:0] Checking_FPU_covSum		//Jaewon_FPU_regstate
);
  assign Checking_FPU_regstate = FPU_state; 	//Jaewon_FPU_regstate
  assign Checking_FPU_covSum = FPU_covSum; 	//Jaewon_FPU_covSum
  wire [31:0] fp_decoder_io_inst; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_wen; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_ren1; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_ren2; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_ren3; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_swap12; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_swap23; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_singleIn; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_singleOut; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_fromint; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_toint; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_fastpipe; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_fma; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_div; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_sqrt; // @[FPU.scala 694:26]
  wire  fp_decoder_io_sigs_wflags; // @[FPU.scala 694:26]
  wire [29:0] fp_decoder_io_covSum; // @[FPU.scala 694:26]
  wire  fp_decoder_metaAssert; // @[FPU.scala 694:26]
  reg [64:0] regfile [0:31]; // @[FPU.scala 748:20]
  reg [95:0] _RAND_0;
  wire [64:0] regfile_ex_rs_0_data; // @[FPU.scala 748:20]
  wire [4:0] regfile_ex_rs_0_addr; // @[FPU.scala 748:20]
  wire [64:0] regfile_ex_rs_1_data; // @[FPU.scala 748:20]
  wire [4:0] regfile_ex_rs_1_addr; // @[FPU.scala 748:20]
  wire [64:0] regfile_ex_rs_2_data; // @[FPU.scala 748:20]
  wire [4:0] regfile_ex_rs_2_addr; // @[FPU.scala 748:20]
  wire [64:0] regfile__T_251_data; // @[FPU.scala 748:20]
  wire [4:0] regfile__T_251_addr; // @[FPU.scala 748:20]
  wire  regfile__T_251_mask; // @[FPU.scala 748:20]
  wire  regfile__T_251_en; // @[FPU.scala 748:20]
  wire [64:0] regfile__T_818_data; // @[FPU.scala 748:20]
  wire [4:0] regfile__T_818_addr; // @[FPU.scala 748:20]
  wire  regfile__T_818_mask; // @[FPU.scala 748:20]
  wire  regfile__T_818_en; // @[FPU.scala 748:20]
  wire  sfma_clock; // @[FPU.scala 795:20]
  wire  sfma_reset; // @[FPU.scala 795:20]
  wire  sfma_io_in_valid; // @[FPU.scala 795:20]
  wire  sfma_io_in_bits_ren3; // @[FPU.scala 795:20]
  wire  sfma_io_in_bits_swap23; // @[FPU.scala 795:20]
  wire [2:0] sfma_io_in_bits_rm; // @[FPU.scala 795:20]
  wire [1:0] sfma_io_in_bits_fmaCmd; // @[FPU.scala 795:20]
  wire [64:0] sfma_io_in_bits_in1; // @[FPU.scala 795:20]
  wire [64:0] sfma_io_in_bits_in2; // @[FPU.scala 795:20]
  wire [64:0] sfma_io_in_bits_in3; // @[FPU.scala 795:20]
  wire [64:0] sfma_io_out_bits_data; // @[FPU.scala 795:20]
  wire [4:0] sfma_io_out_bits_exc; // @[FPU.scala 795:20]
  wire [29:0] sfma_io_covSum; // @[FPU.scala 795:20]
  wire  sfma_metaAssert; // @[FPU.scala 795:20]
  wire  sfma_metaReset; // @[FPU.scala 795:20]
  wire  sfma_fma_halt; // @[FPU.scala 795:20]
  wire  fpiu_clock; // @[FPU.scala 799:20]
  wire  fpiu_io_in_valid; // @[FPU.scala 799:20]
  wire  fpiu_io_in_bits_ren2; // @[FPU.scala 799:20]
  wire  fpiu_io_in_bits_singleIn; // @[FPU.scala 799:20]
  wire  fpiu_io_in_bits_singleOut; // @[FPU.scala 799:20]
  wire  fpiu_io_in_bits_wflags; // @[FPU.scala 799:20]
  wire [2:0] fpiu_io_in_bits_rm; // @[FPU.scala 799:20]
  wire [1:0] fpiu_io_in_bits_typ; // @[FPU.scala 799:20]
  wire [64:0] fpiu_io_in_bits_in1; // @[FPU.scala 799:20]
  wire [64:0] fpiu_io_in_bits_in2; // @[FPU.scala 799:20]
  wire [2:0] fpiu_io_out_bits_in_rm; // @[FPU.scala 799:20]
  wire [64:0] fpiu_io_out_bits_in_in1; // @[FPU.scala 799:20]
  wire [64:0] fpiu_io_out_bits_in_in2; // @[FPU.scala 799:20]
  wire  fpiu_io_out_bits_lt; // @[FPU.scala 799:20]
  wire [63:0] fpiu_io_out_bits_store; // @[FPU.scala 799:20]
  wire [63:0] fpiu_io_out_bits_toint; // @[FPU.scala 799:20]
  wire [4:0] fpiu_io_out_bits_exc; // @[FPU.scala 799:20]
  wire [29:0] fpiu_io_covSum; // @[FPU.scala 799:20]
  wire  fpiu_metaAssert; // @[FPU.scala 799:20]
  wire  fpiu_metaReset; // @[FPU.scala 799:20]
  wire  ifpu_clock; // @[FPU.scala 809:20]
  wire  ifpu_reset; // @[FPU.scala 809:20]
  wire  ifpu_io_in_valid; // @[FPU.scala 809:20]
  wire  ifpu_io_in_bits_singleIn; // @[FPU.scala 809:20]
  wire  ifpu_io_in_bits_wflags; // @[FPU.scala 809:20]
  wire [2:0] ifpu_io_in_bits_rm; // @[FPU.scala 809:20]
  wire [1:0] ifpu_io_in_bits_typ; // @[FPU.scala 809:20]
  wire [63:0] ifpu_io_in_bits_in1; // @[FPU.scala 809:20]
  wire [64:0] ifpu_io_out_bits_data; // @[FPU.scala 809:20]
  wire [4:0] ifpu_io_out_bits_exc; // @[FPU.scala 809:20]
  wire [29:0] ifpu_io_covSum; // @[FPU.scala 809:20]
  wire  ifpu_metaAssert; // @[FPU.scala 809:20]
  wire  ifpu_metaReset; // @[FPU.scala 809:20]
  wire  fpmu_clock; // @[FPU.scala 814:20]
  wire  fpmu_reset; // @[FPU.scala 814:20]
  wire  fpmu_io_in_valid; // @[FPU.scala 814:20]
  wire  fpmu_io_in_bits_ren2; // @[FPU.scala 814:20]
  wire  fpmu_io_in_bits_singleOut; // @[FPU.scala 814:20]
  wire  fpmu_io_in_bits_wflags; // @[FPU.scala 814:20]
  wire [2:0] fpmu_io_in_bits_rm; // @[FPU.scala 814:20]
  wire [64:0] fpmu_io_in_bits_in1; // @[FPU.scala 814:20]
  wire [64:0] fpmu_io_in_bits_in2; // @[FPU.scala 814:20]
  wire [64:0] fpmu_io_out_bits_data; // @[FPU.scala 814:20]
  wire [4:0] fpmu_io_out_bits_exc; // @[FPU.scala 814:20]
  wire  fpmu_io_lt; // @[FPU.scala 814:20]
  wire [29:0] fpmu_io_covSum; // @[FPU.scala 814:20]
  wire  fpmu_metaAssert; // @[FPU.scala 814:20]
  wire  fpmu_metaReset; // @[FPU.scala 814:20]
  wire  dfma_clock; // @[FPU.scala 833:28]
  wire  dfma_reset; // @[FPU.scala 833:28]
  wire  dfma_io_in_valid; // @[FPU.scala 833:28]
  wire  dfma_io_in_bits_ren3; // @[FPU.scala 833:28]
  wire  dfma_io_in_bits_swap23; // @[FPU.scala 833:28]
  wire [2:0] dfma_io_in_bits_rm; // @[FPU.scala 833:28]
  wire [1:0] dfma_io_in_bits_fmaCmd; // @[FPU.scala 833:28]
  wire [64:0] dfma_io_in_bits_in1; // @[FPU.scala 833:28]
  wire [64:0] dfma_io_in_bits_in2; // @[FPU.scala 833:28]
  wire [64:0] dfma_io_in_bits_in3; // @[FPU.scala 833:28]
  wire [64:0] dfma_io_out_bits_data; // @[FPU.scala 833:28]
  wire [4:0] dfma_io_out_bits_exc; // @[FPU.scala 833:28]
  wire [29:0] dfma_io_covSum; // @[FPU.scala 833:28]
  wire  dfma_metaAssert; // @[FPU.scala 833:28]
  wire  dfma_metaReset; // @[FPU.scala 833:28]
  wire  dfma_fma_halt; // @[FPU.scala 833:28]
  wire  divSqrt_clock; // @[FPU.scala 926:27]
  wire  divSqrt_reset; // @[FPU.scala 926:27]
  wire  divSqrt_io_inReady; // @[FPU.scala 926:27]
  wire  divSqrt_io_inValid; // @[FPU.scala 926:27]
  wire  divSqrt_io_sqrtOp; // @[FPU.scala 926:27]
  wire [32:0] divSqrt_io_a; // @[FPU.scala 926:27]
  wire [32:0] divSqrt_io_b; // @[FPU.scala 926:27]
  wire [2:0] divSqrt_io_roundingMode; // @[FPU.scala 926:27]
  wire  divSqrt_io_outValid_div; // @[FPU.scala 926:27]
  wire  divSqrt_io_outValid_sqrt; // @[FPU.scala 926:27]
  wire [32:0] divSqrt_io_out; // @[FPU.scala 926:27]
  wire [4:0] divSqrt_io_exceptionFlags; // @[FPU.scala 926:27]
  wire [29:0] divSqrt_io_covSum; // @[FPU.scala 926:27]
  wire  divSqrt_metaAssert; // @[FPU.scala 926:27]
  wire  divSqrt_metaReset; // @[FPU.scala 926:27]
  wire  divSqrt_divSqrtRecFNToRaw_halt; // @[FPU.scala 926:27]
  wire  divSqrt_1_clock; // @[FPU.scala 926:27]
  wire  divSqrt_1_reset; // @[FPU.scala 926:27]
  wire  divSqrt_1_io_inReady; // @[FPU.scala 926:27]
  wire  divSqrt_1_io_inValid; // @[FPU.scala 926:27]
  wire  divSqrt_1_io_sqrtOp; // @[FPU.scala 926:27]
  wire [64:0] divSqrt_1_io_a; // @[FPU.scala 926:27]
  wire [64:0] divSqrt_1_io_b; // @[FPU.scala 926:27]
  wire [2:0] divSqrt_1_io_roundingMode; // @[FPU.scala 926:27]
  wire  divSqrt_1_io_outValid_div; // @[FPU.scala 926:27]
  wire  divSqrt_1_io_outValid_sqrt; // @[FPU.scala 926:27]
  wire [64:0] divSqrt_1_io_out; // @[FPU.scala 926:27]
  wire [4:0] divSqrt_1_io_exceptionFlags; // @[FPU.scala 926:27]
  wire [29:0] divSqrt_1_io_covSum; // @[FPU.scala 926:27]
  wire  divSqrt_1_metaAssert; // @[FPU.scala 926:27]
  wire  divSqrt_1_metaReset; // @[FPU.scala 926:27]
  wire  divSqrt_1_divSqrtRecFNToRaw_halt; // @[FPU.scala 926:27]
  reg  ex_reg_valid; // @[FPU.scala 698:25]
  reg [31:0] _RAND_1;
  reg [31:0] ex_reg_inst; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg  ex_reg_ctrl_ren2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg  ex_reg_ctrl_ren3; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  ex_reg_ctrl_swap23; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  ex_reg_ctrl_singleIn; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  ex_reg_ctrl_singleOut; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg  ex_reg_ctrl_fromint; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg  ex_reg_ctrl_toint; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg  ex_reg_ctrl_fastpipe; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg  ex_reg_ctrl_fma; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg  ex_reg_ctrl_div; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg  ex_reg_ctrl_sqrt; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg  ex_reg_ctrl_wflags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [4:0] ex_ra_0; // @[FPU.scala 701:31]
  reg [31:0] _RAND_15;
  reg [4:0] ex_ra_1; // @[FPU.scala 701:31]
  reg [31:0] _RAND_16;
  reg [4:0] ex_ra_2; // @[FPU.scala 701:31]
  reg [31:0] _RAND_17;
  reg  load_wb; // @[FPU.scala 704:20]
  reg [31:0] _RAND_18;
  reg  load_wb_double; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [63:0] load_wb_data; // @[Reg.scala 15:16]
  reg [63:0] _RAND_20;
  reg [4:0] load_wb_tag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg  mem_reg_valid; // @[FPU.scala 715:30]
  reg [31:0] _RAND_22;
  wire  killm; // @[FPU.scala 716:25]
  wire  _T_3; // @[FPU.scala 720:41]
  wire  killx; // @[FPU.scala 720:24]
  wire  _T_5; // @[FPU.scala 721:33]
  reg [31:0] mem_reg_inst; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  wire  _T_9; // @[FPU.scala 723:45]
  reg  wb_reg_valid; // @[FPU.scala 723:25]
  reg [31:0] _RAND_24;
  reg  mem_ctrl_singleOut; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg  mem_ctrl_fromint; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg  mem_ctrl_toint; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg  mem_ctrl_fastpipe; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg  mem_ctrl_fma; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg  mem_ctrl_div; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg  mem_ctrl_sqrt; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg  mem_ctrl_wflags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg  wb_ctrl_toint; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  wire [63:0] _T_13; // @[package.scala 32:76]
  wire [63:0] _T_14; // @[FPU.scala 379:23]
  wire  _T_18; // @[rawFloatFromFN.scala 50:34]
  wire  _T_19; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_72; // @[Mux.scala 47:69]
  wire [5:0] _T_73; // @[Mux.scala 47:69]
  wire [5:0] _T_74; // @[Mux.scala 47:69]
  wire [5:0] _T_75; // @[Mux.scala 47:69]
  wire [5:0] _T_76; // @[Mux.scala 47:69]
  wire [5:0] _T_77; // @[Mux.scala 47:69]
  wire [5:0] _T_78; // @[Mux.scala 47:69]
  wire [5:0] _T_79; // @[Mux.scala 47:69]
  wire [5:0] _T_80; // @[Mux.scala 47:69]
  wire [5:0] _T_81; // @[Mux.scala 47:69]
  wire [5:0] _T_82; // @[Mux.scala 47:69]
  wire [5:0] _T_83; // @[Mux.scala 47:69]
  wire [5:0] _T_84; // @[Mux.scala 47:69]
  wire [5:0] _T_85; // @[Mux.scala 47:69]
  wire [5:0] _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_106; // @[Mux.scala 47:69]
  wire [5:0] _T_107; // @[Mux.scala 47:69]
  wire [5:0] _T_108; // @[Mux.scala 47:69]
  wire [5:0] _T_109; // @[Mux.scala 47:69]
  wire [5:0] _T_110; // @[Mux.scala 47:69]
  wire [5:0] _T_111; // @[Mux.scala 47:69]
  wire [5:0] _T_112; // @[Mux.scala 47:69]
  wire [5:0] _T_113; // @[Mux.scala 47:69]
  wire [5:0] _T_114; // @[Mux.scala 47:69]
  wire [5:0] _T_115; // @[Mux.scala 47:69]
  wire [5:0] _T_116; // @[Mux.scala 47:69]
  wire [5:0] _T_117; // @[Mux.scala 47:69]
  wire [5:0] _T_118; // @[Mux.scala 47:69]
  wire [5:0] _T_119; // @[Mux.scala 47:69]
  wire [5:0] _T_120; // @[Mux.scala 47:69]
  wire [5:0] _T_121; // @[Mux.scala 47:69]
  wire [5:0] _T_122; // @[Mux.scala 47:69]
  wire [114:0] _GEN_167; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_123; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_125; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_168; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_126; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_127; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_128; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_169; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_129; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_170; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_131; // @[rawFloatFromFN.scala 59:15]
  wire  _T_132; // @[rawFloatFromFN.scala 62:34]
  wire  _T_134; // @[rawFloatFromFN.scala 63:62]
  wire  _T_137; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_140; // @[rawFloatFromFN.scala 70:48]
  wire [51:0] _T_142; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_144; // @[Cat.scala 29:58]
  wire [2:0] _T_146; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_171; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_148; // @[recFNFromFN.scala 48:79]
  wire [64:0] _T_153; // @[Cat.scala 29:58]
  wire  _T_157; // @[rawFloatFromFN.scala 50:34]
  wire  _T_158; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_182; // @[Mux.scala 47:69]
  wire [4:0] _T_183; // @[Mux.scala 47:69]
  wire [4:0] _T_184; // @[Mux.scala 47:69]
  wire [4:0] _T_185; // @[Mux.scala 47:69]
  wire [4:0] _T_186; // @[Mux.scala 47:69]
  wire [4:0] _T_187; // @[Mux.scala 47:69]
  wire [4:0] _T_188; // @[Mux.scala 47:69]
  wire [4:0] _T_189; // @[Mux.scala 47:69]
  wire [4:0] _T_190; // @[Mux.scala 47:69]
  wire [4:0] _T_191; // @[Mux.scala 47:69]
  wire [4:0] _T_192; // @[Mux.scala 47:69]
  wire [4:0] _T_193; // @[Mux.scala 47:69]
  wire [4:0] _T_194; // @[Mux.scala 47:69]
  wire [4:0] _T_195; // @[Mux.scala 47:69]
  wire [4:0] _T_196; // @[Mux.scala 47:69]
  wire [4:0] _T_197; // @[Mux.scala 47:69]
  wire [4:0] _T_198; // @[Mux.scala 47:69]
  wire [4:0] _T_199; // @[Mux.scala 47:69]
  wire [4:0] _T_200; // @[Mux.scala 47:69]
  wire [4:0] _T_201; // @[Mux.scala 47:69]
  wire [4:0] _T_202; // @[Mux.scala 47:69]
  wire [4:0] _T_203; // @[Mux.scala 47:69]
  wire [53:0] _GEN_172; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_204; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_206; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_173; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_207; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_208; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_209; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_174; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_210; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_175; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_212; // @[rawFloatFromFN.scala 59:15]
  wire  _T_213; // @[rawFloatFromFN.scala 62:34]
  wire  _T_215; // @[rawFloatFromFN.scala 63:62]
  wire  _T_218; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_221; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_223; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_225; // @[Cat.scala 29:58]
  wire [2:0] _T_227; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_176; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_229; // @[recFNFromFN.scala 48:79]
  wire [32:0] _T_234; // @[Cat.scala 29:58]
  wire  _T_237; // @[FPU.scala 286:42]
  wire [64:0] _T_248; // @[Cat.scala 29:58]
  wire  _T_250; // @[FPU.scala 203:56]
  wire [64:0] wdata; // @[FPU.scala 292:8]
  wire  _T_262; // @[FPU.scala 203:56]
  wire  _T_266; // @[FPU.scala 333:96]
  wire  _T_267; // @[FPU.scala 333:55]
  wire  _T_268; // @[FPU.scala 333:31]
  wire  _T_271; // @[FPU.scala 752:11]
  wire  _T_371; // @[FPU.scala 769:29]
  wire  _T_375; // @[FPU.scala 773:38]
  wire  _T_377; // @[FPU.scala 796:33]
  wire  tag; // @[FPU.scala 777:15]
  wire [32:0] _T_383; // @[Cat.scala 29:58]
  wire  _T_385; // @[FPU.scala 280:84]
  wire [32:0] _T_406; // @[FPU.scala 320:31]
  wire [32:0] _T_407; // @[FPU.scala 320:26]
  wire [32:0] _T_412; // @[Cat.scala 29:58]
  wire  _T_414; // @[FPU.scala 280:84]
  wire [32:0] _T_435; // @[FPU.scala 320:31]
  wire [32:0] _T_436; // @[FPU.scala 320:26]
  wire [32:0] _T_441; // @[Cat.scala 29:58]
  wire  _T_443; // @[FPU.scala 280:84]
  wire [32:0] _T_464; // @[FPU.scala 320:31]
  wire [32:0] _T_465; // @[FPU.scala 320:26]
  wire  _T_470; // @[FPU.scala 784:53]
  wire [1:0] _GEN_177; // @[FPU.scala 784:36]
  wire  _T_472; // @[FPU.scala 800:51]
  wire  _T_473; // @[FPU.scala 800:66]
  wire  _T_474; // @[FPU.scala 800:103]
  wire  _T_475; // @[FPU.scala 800:82]
  wire [75:0] _T_485; // @[FPU.scala 231:28]
  wire [11:0] _GEN_178; // @[FPU.scala 234:31]
  wire [11:0] _T_489; // @[FPU.scala 234:31]
  wire [11:0] _T_491; // @[FPU.scala 234:48]
  wire  _T_492; // @[FPU.scala 235:19]
  wire  _T_493; // @[FPU.scala 235:36]
  wire  _T_494; // @[FPU.scala 235:25]
  wire [11:0] _T_496; // @[Cat.scala 29:58]
  wire [11:0] _T_498; // @[FPU.scala 235:10]
  wire [64:0] _T_500; // @[Cat.scala 29:58]
  wire  _T_505; // @[package.scala 32:76]
  wire [64:0] _T_507; // @[package.scala 32:76]
  wire [75:0] _T_517; // @[FPU.scala 231:28]
  wire [11:0] _GEN_179; // @[FPU.scala 234:31]
  wire [11:0] _T_521; // @[FPU.scala 234:31]
  wire [11:0] _T_523; // @[FPU.scala 234:48]
  wire  _T_524; // @[FPU.scala 235:19]
  wire  _T_525; // @[FPU.scala 235:36]
  wire  _T_526; // @[FPU.scala 235:25]
  wire [11:0] _T_528; // @[Cat.scala 29:58]
  wire [11:0] _T_530; // @[FPU.scala 235:10]
  wire [64:0] _T_532; // @[Cat.scala 29:58]
  wire  _T_537; // @[package.scala 32:76]
  wire [64:0] _T_539; // @[package.scala 32:76]
  wire [64:0] _T_582; // @[FPU.scala 812:29]
  reg [4:0] divSqrt_waddr; // @[FPU.scala 821:26]
  reg [31:0] _RAND_34;
  wire  _T_682; // @[FPU.scala 831:56]
  wire [1:0] _T_683; // @[FPU.scala 840:23]
  wire  _T_685; // @[FPU.scala 836:62]
  wire [2:0] _T_686; // @[FPU.scala 840:23]
  wire  _T_687; // @[FPU.scala 840:78]
  wire [1:0] _GEN_186; // @[FPU.scala 840:78]
  wire [1:0] _T_688; // @[FPU.scala 840:78]
  wire [2:0] _GEN_187; // @[FPU.scala 840:78]
  wire [2:0] memLatencyMask; // @[FPU.scala 840:78]
  reg [2:0] wen; // @[FPU.scala 854:16]
  reg [31:0] _RAND_35;
  reg [4:0] wbInfo_0_rd; // @[FPU.scala 855:19]
  reg [31:0] _RAND_36;
  reg  wbInfo_0_single; // @[FPU.scala 855:19]
  reg [31:0] _RAND_37;
  reg [1:0] wbInfo_0_pipeid; // @[FPU.scala 855:19]
  reg [31:0] _RAND_38;
  reg [4:0] wbInfo_1_rd; // @[FPU.scala 855:19]
  reg [31:0] _RAND_39;
  reg  wbInfo_1_single; // @[FPU.scala 855:19]
  reg [31:0] _RAND_40;
  reg [1:0] wbInfo_1_pipeid; // @[FPU.scala 855:19]
  reg [31:0] _RAND_41;
  reg [4:0] wbInfo_2_rd; // @[FPU.scala 855:19]
  reg [31:0] _RAND_42;
  reg  wbInfo_2_single; // @[FPU.scala 855:19]
  reg [31:0] _RAND_43;
  reg [1:0] wbInfo_2_pipeid; // @[FPU.scala 855:19]
  reg [31:0] _RAND_44;
  wire  _T_689; // @[FPU.scala 856:48]
  wire  _T_690; // @[FPU.scala 856:69]
  wire  mem_wen; // @[FPU.scala 856:31]
  wire [1:0] _T_691; // @[FPU.scala 840:23]
  wire [1:0] _T_692; // @[FPU.scala 840:23]
  wire  _T_693; // @[FPU.scala 831:56]
  wire [2:0] _T_694; // @[FPU.scala 840:23]
  wire  _T_696; // @[FPU.scala 836:62]
  wire [3:0] _T_697; // @[FPU.scala 840:23]
  wire [1:0] _T_698; // @[FPU.scala 840:78]
  wire [2:0] _GEN_188; // @[FPU.scala 840:78]
  wire [2:0] _T_699; // @[FPU.scala 840:78]
  wire [3:0] _GEN_189; // @[FPU.scala 840:78]
  wire [3:0] _T_700; // @[FPU.scala 840:78]
  wire [3:0] _GEN_190; // @[FPU.scala 857:62]
  wire [3:0] _T_701; // @[FPU.scala 857:62]
  wire  _T_702; // @[FPU.scala 857:89]
  wire  _T_703; // @[FPU.scala 857:43]
  wire [2:0] _T_704; // @[FPU.scala 840:23]
  wire [2:0] _T_705; // @[FPU.scala 840:23]
  wire [3:0] _T_707; // @[FPU.scala 840:23]
  wire [4:0] _T_710; // @[FPU.scala 840:23]
  wire [2:0] _T_711; // @[FPU.scala 840:78]
  wire [3:0] _GEN_191; // @[FPU.scala 840:78]
  wire [3:0] _T_712; // @[FPU.scala 840:78]
  wire [4:0] _GEN_192; // @[FPU.scala 840:78]
  wire [4:0] _T_713; // @[FPU.scala 840:78]
  wire [4:0] _GEN_193; // @[FPU.scala 857:101]
  wire [4:0] _T_714; // @[FPU.scala 857:101]
  wire  _T_715; // @[FPU.scala 857:128]
  wire  _T_716; // @[FPU.scala 857:93]
  reg  write_port_busy; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  wire [2:0] _GEN_194; // @[FPU.scala 866:23]
  wire [2:0] _T_723; // @[FPU.scala 866:23]
  wire  _T_726; // @[FPU.scala 869:30]
  wire [1:0] _T_733; // @[FPU.scala 842:63]
  wire [1:0] _GEN_195; // @[FPU.scala 842:108]
  wire [1:0] _T_735; // @[FPU.scala 842:108]
  wire [1:0] _T_736; // @[FPU.scala 842:108]
  wire  _T_740; // @[FPU.scala 869:30]
  wire  _T_754; // @[FPU.scala 869:30]
  wire  divSqrt_typeTag; // @[FPU.scala 941:37]
  reg  divSqrt_killed; // @[FPU.scala 919:29]
  reg [31:0] _RAND_46;
  wire  _T_1007; // @[FPU.scala 941:37]
  wire  _GEN_156; // @[FPU.scala 941:66]
  wire  divSqrt_wen; // @[FPU.scala 941:66]
  wire  wdouble; // @[FPU.scala 879:20]
  wire  _T_767; // @[package.scala 32:86]
  wire [64:0] _T_768; // @[package.scala 32:76]
  wire  _T_769; // @[package.scala 32:86]
  wire [64:0] _T_770; // @[package.scala 32:76]
  wire  _T_771; // @[package.scala 32:86]
  wire [64:0] _T_772; // @[package.scala 32:76]
  wire  _T_1023; // @[FPU.scala 203:56]
  wire [64:0] _T_1021; // @[FPU.scala 361:25]
  wire [64:0] _T_1024; // @[FPU.scala 362:10]
  wire [32:0] _GEN_157; // @[FPU.scala 941:66]
  wire [64:0] divSqrt_wdata; // @[FPU.scala 941:66]
  wire [64:0] _T_773; // @[FPU.scala 880:22]
  wire  _T_774; // @[FPU.scala 286:42]
  wire [64:0] _T_783; // @[Cat.scala 29:58]
  wire  _T_784; // @[FPU.scala 203:56]
  wire [64:0] _T_785; // @[FPU.scala 292:8]
  wire [64:0] wdata_1; // @[package.scala 32:76]
  wire [4:0] _T_789; // @[package.scala 32:76]
  wire [4:0] _T_791; // @[package.scala 32:76]
  wire [4:0] wexc; // @[package.scala 32:76]
  wire  frfWriteBundle_1_wrenf; // @[FPU.scala 882:35]
  wire  _T_807; // @[FPU.scala 203:56]
  wire  _T_811; // @[FPU.scala 333:96]
  wire  _T_812; // @[FPU.scala 333:55]
  wire  _T_813; // @[FPU.scala 333:31]
  wire  _T_816; // @[FPU.scala 883:11]
  wire  wb_toint_valid; // @[FPU.scala 898:37]
  reg [4:0] wb_toint_exc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  wire  _T_907; // @[FPU.scala 900:41]
  wire [4:0] _T_910; // @[FPU.scala 902:8]
  wire [4:0] _GEN_158; // @[FPU.scala 941:66]
  wire [4:0] divSqrt_flags; // @[FPU.scala 941:66]
  wire [4:0] _T_911; // @[FPU.scala 903:8]
  wire [4:0] _T_912; // @[FPU.scala 902:48]
  wire [4:0] _T_914; // @[FPU.scala 904:8]
  wire  _T_916; // @[FPU.scala 906:47]
  wire  _T_917; // @[FPU.scala 906:72]
  wire  divSqrt_write_port_busy; // @[FPU.scala 906:65]
  wire  _T_918; // @[FPU.scala 907:33]
  wire  _T_919; // @[FPU.scala 907:68]
  wire  _T_920; // @[FPU.scala 907:51]
  wire  _T_922; // @[FPU.scala 907:87]
  wire  _T_924; // @[FPU.scala 907:120]
  wire  divSqrt_inFlight; // @[FPU.scala 934:34]
  wire  _T_925; // @[FPU.scala 907:131]
  wire  _T_927; // @[FPU.scala 908:34]
  wire  _T_934; // @[FPU.scala 911:96]
  reg  _T_936; // @[FPU.scala 911:55]
  reg [31:0] _RAND_48;
  wire  _T_942; // @[FPU.scala 912:60]
  wire  _T_947; // @[package.scala 15:47]
  wire  _T_948; // @[package.scala 15:47]
  wire  _T_949; // @[package.scala 64:59]
  wire  _T_951; // @[FPU.scala 916:67]
  wire  _T_952; // @[FPU.scala 916:87]
  wire  _T_953; // @[FPU.scala 916:73]
  wire  _T_961; // @[FPU.scala 927:43]
  wire  _T_963; // @[FPU.scala 927:65]
  wire [75:0] _T_969; // @[FPU.scala 231:28]
  wire [11:0] _T_973; // @[FPU.scala 234:31]
  wire [11:0] _T_975; // @[FPU.scala 234:48]
  wire  _T_976; // @[FPU.scala 235:19]
  wire  _T_977; // @[FPU.scala 235:36]
  wire  _T_978; // @[FPU.scala 235:25]
  wire [8:0] _T_980; // @[Cat.scala 29:58]
  wire [8:0] _T_982; // @[FPU.scala 235:10]
  wire [9:0] _T_983; // @[Cat.scala 29:58]
  wire [75:0] _T_988; // @[FPU.scala 231:28]
  wire [11:0] _T_992; // @[FPU.scala 234:31]
  wire [11:0] _T_994; // @[FPU.scala 234:48]
  wire  _T_995; // @[FPU.scala 235:19]
  wire  _T_996; // @[FPU.scala 235:36]
  wire  _T_997; // @[FPU.scala 235:25]
  wire [8:0] _T_999; // @[Cat.scala 29:58]
  wire [8:0] _T_1001; // @[FPU.scala 235:10]
  wire [9:0] _T_1002; // @[Cat.scala 29:58]
  wire  _T_1005; // @[FPU.scala 936:32]
  wire  _T_1010; // @[FPU.scala 927:43]
  wire  _T_1012; // @[FPU.scala 927:65]
  wire  _T_1016; // @[FPU.scala 936:32]
  reg [19:0] FPU_state; // @[Register tracking FPU state]
  reg [31:0] _RAND_49;
  reg  FPU_cov [0:1048575]; // @[Coverage map for FPU]
  reg [31:0] _RAND_50;
  wire  FPU_cov_read_data; // @[Coverage map for FPU]
  wire [19:0] FPU_cov_read_addr; // @[Coverage map for FPU]
  wire  FPU_cov_write_data; // @[Coverage map for FPU]
  wire [19:0] FPU_cov_write_addr; // @[Coverage map for FPU]
  wire  FPU_cov_write_mask; // @[Coverage map for FPU]
  wire  FPU_cov_write_en; // @[Coverage map for FPU]
  reg [29:0] FPU_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_51;
  wire  wbInfo_0_single_shl;
  wire [19:0] wbInfo_0_single_pad;
  wire [16:0] ex_reg_ctrl_fromint_shl;
  wire [19:0] ex_reg_ctrl_fromint_pad;
  wire [19:0] wb_ctrl_toint_shl;
  wire [19:0] wb_ctrl_toint_pad;
  wire [13:0] ex_reg_ctrl_fastpipe_shl;
  wire [19:0] ex_reg_ctrl_fastpipe_pad;
  wire [1:0] mem_reg_valid_shl;
  wire [19:0] mem_reg_valid_pad;
  wire [14:0] write_port_busy_shl;
  wire [19:0] write_port_busy_pad;
  wire [2:0] ex_reg_ctrl_singleIn_shl;
  wire [19:0] ex_reg_ctrl_singleIn_pad;
  wire [1:0] mem_ctrl_fastpipe_shl;
  wire [19:0] mem_ctrl_fastpipe_pad;
  wire [13:0] wbInfo_0_pipeid_shl;
  wire [19:0] wbInfo_0_pipeid_pad;
  wire [1:0] load_wb_double_shl;
  wire [19:0] load_wb_double_pad;
  wire  ex_reg_ctrl_singleOut_shl;
  wire [19:0] ex_reg_ctrl_singleOut_pad;
  wire [3:0] wen_shl;
  wire [19:0] wen_pad;
  wire [14:0] mem_ctrl_toint_shl;
  wire [19:0] mem_ctrl_toint_pad;
  wire [7:0] wb_reg_valid_shl;
  wire [19:0] wb_reg_valid_pad;
  wire [2:0] ex_reg_ctrl_fma_shl;
  wire [19:0] ex_reg_ctrl_fma_pad;
  wire [4:0] mem_ctrl_singleOut_shl;
  wire [19:0] mem_ctrl_singleOut_pad;
  wire [8:0] mem_ctrl_fromint_shl;
  wire [19:0] mem_ctrl_fromint_pad;
  wire [17:0] mem_ctrl_fma_shl;
  wire [19:0] mem_ctrl_fma_pad;
  wire [7:0] ex_reg_valid_shl;
  wire [19:0] ex_reg_valid_pad;
  wire [16:0] divSqrt_killed_shl;
  wire [19:0] divSqrt_killed_pad;
  wire [19:0] FPU_xor7;
  wire [19:0] FPU_xor18;
  wire [19:0] FPU_xor8;
  wire [19:0] FPU_xor3;
  wire [19:0] FPU_xor9;
  wire [19:0] FPU_xor22;
  wire [19:0] FPU_xor10;
  wire [19:0] FPU_xor4;
  wire [19:0] FPU_xor1;
  wire [19:0] FPU_xor11;
  wire [19:0] FPU_xor26;
  wire [19:0] FPU_xor12;
  wire [19:0] FPU_xor5;
  wire [19:0] FPU_xor13;
  wire [19:0] FPU_xor30;
  wire [19:0] FPU_xor14;
  wire [19:0] FPU_xor6;
  wire [19:0] FPU_xor2;
  wire [19:0] FPU_xor0;
  wire [29:0] divSqrt_1_sum;
  wire [29:0] ifpu_sum;
  wire [29:0] divSqrt_sum;
  wire [29:0] fpmu_sum;
  wire [29:0] fp_decoder_sum;
  wire [29:0] dfma_sum;
  wire [29:0] fpiu_sum;
  wire [29:0] sfma_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  ifpu_metaAssert_wire;
  wire  fpmu_metaAssert_wire;
  wire  fp_decoder_metaAssert_wire;
  wire  fpiu_metaAssert_wire;
  wire  divSqrt_1_metaAssert_wire;
  wire  divSqrt_metaAssert_wire;
  wire  dfma_metaAssert_wire;
  wire  sfma_metaAssert_wire;
  wire  FPU_or3;
  wire  FPU_or10;
  wire  FPU_or4;
  wire  FPU_or1;
  wire  FPU_or5;
  wire  FPU_or14;
  wire  FPU_or6;
  wire  FPU_or2;
  wire  FPU_or0;
  reg  FPU_metaAssert;
  reg [31:0] _RAND_52;
  FPUDecoder fp_decoder ( // @[FPU.scala 694:26]
    .io_inst(fp_decoder_io_inst),
    .io_sigs_wen(fp_decoder_io_sigs_wen),
    .io_sigs_ren1(fp_decoder_io_sigs_ren1),
    .io_sigs_ren2(fp_decoder_io_sigs_ren2),
    .io_sigs_ren3(fp_decoder_io_sigs_ren3),
    .io_sigs_swap12(fp_decoder_io_sigs_swap12),
    .io_sigs_swap23(fp_decoder_io_sigs_swap23),
    .io_sigs_singleIn(fp_decoder_io_sigs_singleIn),
    .io_sigs_singleOut(fp_decoder_io_sigs_singleOut),
    .io_sigs_fromint(fp_decoder_io_sigs_fromint),
    .io_sigs_toint(fp_decoder_io_sigs_toint),
    .io_sigs_fastpipe(fp_decoder_io_sigs_fastpipe),
    .io_sigs_fma(fp_decoder_io_sigs_fma),
    .io_sigs_div(fp_decoder_io_sigs_div),
    .io_sigs_sqrt(fp_decoder_io_sigs_sqrt),
    .io_sigs_wflags(fp_decoder_io_sigs_wflags),
    .io_covSum(fp_decoder_io_covSum),
    .metaAssert(fp_decoder_metaAssert)
  );
  FPUFMAPipe sfma ( // @[FPU.scala 795:20]
    .clock(sfma_clock),
    .reset(sfma_reset),
    .io_in_valid(sfma_io_in_valid),
    .io_in_bits_ren3(sfma_io_in_bits_ren3),
    .io_in_bits_swap23(sfma_io_in_bits_swap23),
    .io_in_bits_rm(sfma_io_in_bits_rm),
    .io_in_bits_fmaCmd(sfma_io_in_bits_fmaCmd),
    .io_in_bits_in1(sfma_io_in_bits_in1),
    .io_in_bits_in2(sfma_io_in_bits_in2),
    .io_in_bits_in3(sfma_io_in_bits_in3),
    .io_out_bits_data(sfma_io_out_bits_data),
    .io_out_bits_exc(sfma_io_out_bits_exc),
    .io_covSum(sfma_io_covSum),
    .metaAssert(sfma_metaAssert),
    .metaReset(sfma_metaReset),
    .fma_halt(sfma_fma_halt)
  );
  FPToInt fpiu ( // @[FPU.scala 799:20]
    .clock(fpiu_clock),
    .io_in_valid(fpiu_io_in_valid),
    .io_in_bits_ren2(fpiu_io_in_bits_ren2),
    .io_in_bits_singleIn(fpiu_io_in_bits_singleIn),
    .io_in_bits_singleOut(fpiu_io_in_bits_singleOut),
    .io_in_bits_wflags(fpiu_io_in_bits_wflags),
    .io_in_bits_rm(fpiu_io_in_bits_rm),
    .io_in_bits_typ(fpiu_io_in_bits_typ),
    .io_in_bits_in1(fpiu_io_in_bits_in1),
    .io_in_bits_in2(fpiu_io_in_bits_in2),
    .io_out_bits_in_rm(fpiu_io_out_bits_in_rm),
    .io_out_bits_in_in1(fpiu_io_out_bits_in_in1),
    .io_out_bits_in_in2(fpiu_io_out_bits_in_in2),
    .io_out_bits_lt(fpiu_io_out_bits_lt),
    .io_out_bits_store(fpiu_io_out_bits_store),
    .io_out_bits_toint(fpiu_io_out_bits_toint),
    .io_out_bits_exc(fpiu_io_out_bits_exc),
    .io_covSum(fpiu_io_covSum),
    .metaAssert(fpiu_metaAssert),
    .metaReset(fpiu_metaReset)
  );
  IntToFP ifpu ( // @[FPU.scala 809:20]
    .clock(ifpu_clock),
    .reset(ifpu_reset),
    .io_in_valid(ifpu_io_in_valid),
    .io_in_bits_singleIn(ifpu_io_in_bits_singleIn),
    .io_in_bits_wflags(ifpu_io_in_bits_wflags),
    .io_in_bits_rm(ifpu_io_in_bits_rm),
    .io_in_bits_typ(ifpu_io_in_bits_typ),
    .io_in_bits_in1(ifpu_io_in_bits_in1),
    .io_out_bits_data(ifpu_io_out_bits_data),
    .io_out_bits_exc(ifpu_io_out_bits_exc),
    .io_covSum(ifpu_io_covSum),
    .metaAssert(ifpu_metaAssert),
    .metaReset(ifpu_metaReset)
  );
  FPToFP fpmu ( // @[FPU.scala 814:20]
    .clock(fpmu_clock),
    .reset(fpmu_reset),
    .io_in_valid(fpmu_io_in_valid),
    .io_in_bits_ren2(fpmu_io_in_bits_ren2),
    .io_in_bits_singleOut(fpmu_io_in_bits_singleOut),
    .io_in_bits_wflags(fpmu_io_in_bits_wflags),
    .io_in_bits_rm(fpmu_io_in_bits_rm),
    .io_in_bits_in1(fpmu_io_in_bits_in1),
    .io_in_bits_in2(fpmu_io_in_bits_in2),
    .io_out_bits_data(fpmu_io_out_bits_data),
    .io_out_bits_exc(fpmu_io_out_bits_exc),
    .io_lt(fpmu_io_lt),
    .io_covSum(fpmu_io_covSum),
    .metaAssert(fpmu_metaAssert),
    .metaReset(fpmu_metaReset)
  );
  FPUFMAPipe_1 dfma ( // @[FPU.scala 833:28]
    .clock(dfma_clock),
    .reset(dfma_reset),
    .io_in_valid(dfma_io_in_valid),
    .io_in_bits_ren3(dfma_io_in_bits_ren3),
    .io_in_bits_swap23(dfma_io_in_bits_swap23),
    .io_in_bits_rm(dfma_io_in_bits_rm),
    .io_in_bits_fmaCmd(dfma_io_in_bits_fmaCmd),
    .io_in_bits_in1(dfma_io_in_bits_in1),
    .io_in_bits_in2(dfma_io_in_bits_in2),
    .io_in_bits_in3(dfma_io_in_bits_in3),
    .io_out_bits_data(dfma_io_out_bits_data),
    .io_out_bits_exc(dfma_io_out_bits_exc),
    .io_covSum(dfma_io_covSum),
    .metaAssert(dfma_metaAssert),
    .metaReset(dfma_metaReset),
    .fma_halt(dfma_fma_halt)
  );
  DivSqrtRecFN_small divSqrt ( // @[FPU.scala 926:27]
    .clock(divSqrt_clock),
    .reset(divSqrt_reset),
    .io_inReady(divSqrt_io_inReady),
    .io_inValid(divSqrt_io_inValid),
    .io_sqrtOp(divSqrt_io_sqrtOp),
    .io_a(divSqrt_io_a),
    .io_b(divSqrt_io_b),
    .io_roundingMode(divSqrt_io_roundingMode),
    .io_outValid_div(divSqrt_io_outValid_div),
    .io_outValid_sqrt(divSqrt_io_outValid_sqrt),
    .io_out(divSqrt_io_out),
    .io_exceptionFlags(divSqrt_io_exceptionFlags),
    .io_covSum(divSqrt_io_covSum),
    .metaAssert(divSqrt_metaAssert),
    .metaReset(divSqrt_metaReset),
    .divSqrtRecFNToRaw_halt(divSqrt_divSqrtRecFNToRaw_halt)
  );
  DivSqrtRecFN_small_1 divSqrt_1 ( // @[FPU.scala 926:27]
    .clock(divSqrt_1_clock),
    .reset(divSqrt_1_reset),
    .io_inReady(divSqrt_1_io_inReady),
    .io_inValid(divSqrt_1_io_inValid),
    .io_sqrtOp(divSqrt_1_io_sqrtOp),
    .io_a(divSqrt_1_io_a),
    .io_b(divSqrt_1_io_b),
    .io_roundingMode(divSqrt_1_io_roundingMode),
    .io_outValid_div(divSqrt_1_io_outValid_div),
    .io_outValid_sqrt(divSqrt_1_io_outValid_sqrt),
    .io_out(divSqrt_1_io_out),
    .io_exceptionFlags(divSqrt_1_io_exceptionFlags),
    .io_covSum(divSqrt_1_io_covSum),
    .metaAssert(divSqrt_1_metaAssert),
    .metaReset(divSqrt_1_metaReset),
    .divSqrtRecFNToRaw_halt(divSqrt_1_divSqrtRecFNToRaw_halt)
  );
  assign regfile_ex_rs_0_addr = ex_ra_0;
  assign regfile_ex_rs_0_data = regfile[regfile_ex_rs_0_addr]; // @[FPU.scala 748:20]
  assign regfile_ex_rs_1_addr = ex_ra_1;
  assign regfile_ex_rs_1_data = regfile[regfile_ex_rs_1_addr]; // @[FPU.scala 748:20]
  assign regfile_ex_rs_2_addr = ex_ra_2;
  assign regfile_ex_rs_2_data = regfile[regfile_ex_rs_2_addr]; // @[FPU.scala 748:20]
  assign regfile__T_251_data = _T_250 ? _T_248 : _T_153;
  assign regfile__T_251_addr = load_wb_tag;
  assign regfile__T_251_mask = 1'h1;
  assign regfile__T_251_en = load_wb;
  assign regfile__T_818_data = wdouble ? _T_773 : _T_785;
  assign regfile__T_818_addr = divSqrt_wen ? divSqrt_waddr : wbInfo_0_rd;
  assign regfile__T_818_mask = 1'h1;
  assign regfile__T_818_en = wen[0] | divSqrt_wen;
  assign killm = io_killm | io_nack_mem; // @[FPU.scala 716:25]
  assign _T_3 = mem_reg_valid & killm; // @[FPU.scala 720:41]
  assign killx = io_killx | _T_3; // @[FPU.scala 720:24]
  assign _T_5 = ex_reg_valid & ~killx; // @[FPU.scala 721:33]
  assign _T_9 = mem_reg_valid & ~killm; // @[FPU.scala 723:45]
  assign _T_13 = load_wb_double ? 64'h0 : 64'hffffffff00000000; // @[package.scala 32:76]
  assign _T_14 = _T_13 | load_wb_data; // @[FPU.scala 379:23]
  assign _T_18 = _T_14[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_19 = _T_14[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_72 = _T_14[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  assign _T_73 = _T_14[2] ? 6'h31 : _T_72; // @[Mux.scala 47:69]
  assign _T_74 = _T_14[3] ? 6'h30 : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = _T_14[4] ? 6'h2f : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = _T_14[5] ? 6'h2e : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = _T_14[6] ? 6'h2d : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = _T_14[7] ? 6'h2c : _T_77; // @[Mux.scala 47:69]
  assign _T_79 = _T_14[8] ? 6'h2b : _T_78; // @[Mux.scala 47:69]
  assign _T_80 = _T_14[9] ? 6'h2a : _T_79; // @[Mux.scala 47:69]
  assign _T_81 = _T_14[10] ? 6'h29 : _T_80; // @[Mux.scala 47:69]
  assign _T_82 = _T_14[11] ? 6'h28 : _T_81; // @[Mux.scala 47:69]
  assign _T_83 = _T_14[12] ? 6'h27 : _T_82; // @[Mux.scala 47:69]
  assign _T_84 = _T_14[13] ? 6'h26 : _T_83; // @[Mux.scala 47:69]
  assign _T_85 = _T_14[14] ? 6'h25 : _T_84; // @[Mux.scala 47:69]
  assign _T_86 = _T_14[15] ? 6'h24 : _T_85; // @[Mux.scala 47:69]
  assign _T_87 = _T_14[16] ? 6'h23 : _T_86; // @[Mux.scala 47:69]
  assign _T_88 = _T_14[17] ? 6'h22 : _T_87; // @[Mux.scala 47:69]
  assign _T_89 = _T_14[18] ? 6'h21 : _T_88; // @[Mux.scala 47:69]
  assign _T_90 = _T_14[19] ? 6'h20 : _T_89; // @[Mux.scala 47:69]
  assign _T_91 = _T_14[20] ? 6'h1f : _T_90; // @[Mux.scala 47:69]
  assign _T_92 = _T_14[21] ? 6'h1e : _T_91; // @[Mux.scala 47:69]
  assign _T_93 = _T_14[22] ? 6'h1d : _T_92; // @[Mux.scala 47:69]
  assign _T_94 = _T_14[23] ? 6'h1c : _T_93; // @[Mux.scala 47:69]
  assign _T_95 = _T_14[24] ? 6'h1b : _T_94; // @[Mux.scala 47:69]
  assign _T_96 = _T_14[25] ? 6'h1a : _T_95; // @[Mux.scala 47:69]
  assign _T_97 = _T_14[26] ? 6'h19 : _T_96; // @[Mux.scala 47:69]
  assign _T_98 = _T_14[27] ? 6'h18 : _T_97; // @[Mux.scala 47:69]
  assign _T_99 = _T_14[28] ? 6'h17 : _T_98; // @[Mux.scala 47:69]
  assign _T_100 = _T_14[29] ? 6'h16 : _T_99; // @[Mux.scala 47:69]
  assign _T_101 = _T_14[30] ? 6'h15 : _T_100; // @[Mux.scala 47:69]
  assign _T_102 = _T_14[31] ? 6'h14 : _T_101; // @[Mux.scala 47:69]
  assign _T_103 = _T_14[32] ? 6'h13 : _T_102; // @[Mux.scala 47:69]
  assign _T_104 = _T_14[33] ? 6'h12 : _T_103; // @[Mux.scala 47:69]
  assign _T_105 = _T_14[34] ? 6'h11 : _T_104; // @[Mux.scala 47:69]
  assign _T_106 = _T_14[35] ? 6'h10 : _T_105; // @[Mux.scala 47:69]
  assign _T_107 = _T_14[36] ? 6'hf : _T_106; // @[Mux.scala 47:69]
  assign _T_108 = _T_14[37] ? 6'he : _T_107; // @[Mux.scala 47:69]
  assign _T_109 = _T_14[38] ? 6'hd : _T_108; // @[Mux.scala 47:69]
  assign _T_110 = _T_14[39] ? 6'hc : _T_109; // @[Mux.scala 47:69]
  assign _T_111 = _T_14[40] ? 6'hb : _T_110; // @[Mux.scala 47:69]
  assign _T_112 = _T_14[41] ? 6'ha : _T_111; // @[Mux.scala 47:69]
  assign _T_113 = _T_14[42] ? 6'h9 : _T_112; // @[Mux.scala 47:69]
  assign _T_114 = _T_14[43] ? 6'h8 : _T_113; // @[Mux.scala 47:69]
  assign _T_115 = _T_14[44] ? 6'h7 : _T_114; // @[Mux.scala 47:69]
  assign _T_116 = _T_14[45] ? 6'h6 : _T_115; // @[Mux.scala 47:69]
  assign _T_117 = _T_14[46] ? 6'h5 : _T_116; // @[Mux.scala 47:69]
  assign _T_118 = _T_14[47] ? 6'h4 : _T_117; // @[Mux.scala 47:69]
  assign _T_119 = _T_14[48] ? 6'h3 : _T_118; // @[Mux.scala 47:69]
  assign _T_120 = _T_14[49] ? 6'h2 : _T_119; // @[Mux.scala 47:69]
  assign _T_121 = _T_14[50] ? 6'h1 : _T_120; // @[Mux.scala 47:69]
  assign _T_122 = _T_14[51] ? 6'h0 : _T_121; // @[Mux.scala 47:69]
  assign _GEN_167 = {{63'd0}, _T_14[51:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_123 = _GEN_167 << _T_122; // @[rawFloatFromFN.scala 54:36]
  assign _T_125 = {_T_123[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_168 = {{6'd0}, _T_122}; // @[rawFloatFromFN.scala 57:26]
  assign _T_126 = _GEN_168 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _T_127 = _T_18 ? _T_126 : {{1'd0}, _T_14[62:52]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_128 = _T_18 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_169 = {{9'd0}, _T_128}; // @[rawFloatFromFN.scala 60:22]
  assign _T_129 = 11'h400 | _GEN_169; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_170 = {{1'd0}, _T_129}; // @[rawFloatFromFN.scala 59:15]
  assign _T_131 = _T_127 + _GEN_170; // @[rawFloatFromFN.scala 59:15]
  assign _T_132 = _T_18 & _T_19; // @[rawFloatFromFN.scala 62:34]
  assign _T_134 = _T_131[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_137 = _T_134 & ~_T_19; // @[rawFloatFromFN.scala 66:33]
  assign _T_140 = {1'b0,$signed(_T_131)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_142 = _T_18 ? _T_125 : _T_14[51:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_144 = {1'h0,~_T_132,_T_142}; // @[Cat.scala 29:58]
  assign _T_146 = _T_132 ? 3'h0 : _T_140[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_171 = {{2'd0}, _T_137}; // @[recFNFromFN.scala 48:79]
  assign _T_148 = _T_146 | _GEN_171; // @[recFNFromFN.scala 48:79]
  assign _T_153 = {_T_14[63],_T_148,_T_140[8:0],_T_144[51:0]}; // @[Cat.scala 29:58]
  assign _T_157 = _T_14[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_158 = _T_14[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_182 = _T_14[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _T_183 = _T_14[2] ? 5'h14 : _T_182; // @[Mux.scala 47:69]
  assign _T_184 = _T_14[3] ? 5'h13 : _T_183; // @[Mux.scala 47:69]
  assign _T_185 = _T_14[4] ? 5'h12 : _T_184; // @[Mux.scala 47:69]
  assign _T_186 = _T_14[5] ? 5'h11 : _T_185; // @[Mux.scala 47:69]
  assign _T_187 = _T_14[6] ? 5'h10 : _T_186; // @[Mux.scala 47:69]
  assign _T_188 = _T_14[7] ? 5'hf : _T_187; // @[Mux.scala 47:69]
  assign _T_189 = _T_14[8] ? 5'he : _T_188; // @[Mux.scala 47:69]
  assign _T_190 = _T_14[9] ? 5'hd : _T_189; // @[Mux.scala 47:69]
  assign _T_191 = _T_14[10] ? 5'hc : _T_190; // @[Mux.scala 47:69]
  assign _T_192 = _T_14[11] ? 5'hb : _T_191; // @[Mux.scala 47:69]
  assign _T_193 = _T_14[12] ? 5'ha : _T_192; // @[Mux.scala 47:69]
  assign _T_194 = _T_14[13] ? 5'h9 : _T_193; // @[Mux.scala 47:69]
  assign _T_195 = _T_14[14] ? 5'h8 : _T_194; // @[Mux.scala 47:69]
  assign _T_196 = _T_14[15] ? 5'h7 : _T_195; // @[Mux.scala 47:69]
  assign _T_197 = _T_14[16] ? 5'h6 : _T_196; // @[Mux.scala 47:69]
  assign _T_198 = _T_14[17] ? 5'h5 : _T_197; // @[Mux.scala 47:69]
  assign _T_199 = _T_14[18] ? 5'h4 : _T_198; // @[Mux.scala 47:69]
  assign _T_200 = _T_14[19] ? 5'h3 : _T_199; // @[Mux.scala 47:69]
  assign _T_201 = _T_14[20] ? 5'h2 : _T_200; // @[Mux.scala 47:69]
  assign _T_202 = _T_14[21] ? 5'h1 : _T_201; // @[Mux.scala 47:69]
  assign _T_203 = _T_14[22] ? 5'h0 : _T_202; // @[Mux.scala 47:69]
  assign _GEN_172 = {{31'd0}, _T_14[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_204 = _GEN_172 << _T_203; // @[rawFloatFromFN.scala 54:36]
  assign _T_206 = {_T_204[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_173 = {{4'd0}, _T_203}; // @[rawFloatFromFN.scala 57:26]
  assign _T_207 = _GEN_173 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_208 = _T_157 ? _T_207 : {{1'd0}, _T_14[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_209 = _T_157 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_174 = {{6'd0}, _T_209}; // @[rawFloatFromFN.scala 60:22]
  assign _T_210 = 8'h80 | _GEN_174; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_175 = {{1'd0}, _T_210}; // @[rawFloatFromFN.scala 59:15]
  assign _T_212 = _T_208 + _GEN_175; // @[rawFloatFromFN.scala 59:15]
  assign _T_213 = _T_157 & _T_158; // @[rawFloatFromFN.scala 62:34]
  assign _T_215 = _T_212[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_218 = _T_215 & ~_T_158; // @[rawFloatFromFN.scala 66:33]
  assign _T_221 = {1'b0,$signed(_T_212)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_223 = _T_157 ? _T_206 : _T_14[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_225 = {1'h0,~_T_213,_T_223}; // @[Cat.scala 29:58]
  assign _T_227 = _T_213 ? 3'h0 : _T_221[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_176 = {{2'd0}, _T_218}; // @[recFNFromFN.scala 48:79]
  assign _T_229 = _T_227 | _GEN_176; // @[recFNFromFN.scala 48:79]
  assign _T_234 = {_T_14[31],_T_229,_T_221[5:0],_T_225[22:0]}; // @[Cat.scala 29:58]
  assign _T_237 = &_T_153[51:32]; // @[FPU.scala 286:42]
  assign _T_248 = {_T_153[64:61],_T_237,_T_153[59:53],_T_234[31],_T_153[51:32],_T_234[32],_T_234[30:0]}; // @[Cat.scala 29:58]
  assign _T_250 = &_T_153[63:61]; // @[FPU.scala 203:56]
  assign wdata = _T_250 ? _T_248 : _T_153; // @[FPU.scala 292:8]
  assign _T_262 = &wdata[63:61]; // @[FPU.scala 203:56]
  assign _T_266 = &wdata[51:32]; // @[FPU.scala 333:96]
  assign _T_267 = wdata[60] == _T_266; // @[FPU.scala 333:55]
  assign _T_268 = ~_T_262 | _T_267; // @[FPU.scala 333:31]
  assign _T_271 = _T_268 | reset; // @[FPU.scala 752:11]
  assign _T_371 = ~fp_decoder_io_sigs_swap12 & ~fp_decoder_io_sigs_swap23; // @[FPU.scala 769:29]
  assign _T_375 = ex_reg_inst[14:12] == 3'h7; // @[FPU.scala 773:38]
  assign _T_377 = ex_reg_valid & ex_reg_ctrl_fma; // @[FPU.scala 796:33]
  assign tag = ~ex_reg_ctrl_singleIn; // @[FPU.scala 777:15]
  assign _T_383 = {regfile_ex_rs_0_data[31],regfile_ex_rs_0_data[52],regfile_ex_rs_0_data[30:0]}; // @[Cat.scala 29:58]
  assign _T_385 = &regfile_ex_rs_0_data[64:60]; // @[FPU.scala 280:84]
  assign _T_406 = _T_385 ? 33'h0 : 33'he0400000; // @[FPU.scala 320:31]
  assign _T_407 = _T_383 | _T_406; // @[FPU.scala 320:26]
  assign _T_412 = {regfile_ex_rs_1_data[31],regfile_ex_rs_1_data[52],regfile_ex_rs_1_data[30:0]}; // @[Cat.scala 29:58]
  assign _T_414 = &regfile_ex_rs_1_data[64:60]; // @[FPU.scala 280:84]
  assign _T_435 = _T_414 ? 33'h0 : 33'he0400000; // @[FPU.scala 320:31]
  assign _T_436 = _T_412 | _T_435; // @[FPU.scala 320:26]
  assign _T_441 = {regfile_ex_rs_2_data[31],regfile_ex_rs_2_data[52],regfile_ex_rs_2_data[30:0]}; // @[Cat.scala 29:58]
  assign _T_443 = &regfile_ex_rs_2_data[64:60]; // @[FPU.scala 280:84]
  assign _T_464 = _T_443 ? 33'h0 : 33'he0400000; // @[FPU.scala 320:31]
  assign _T_465 = _T_441 | _T_464; // @[FPU.scala 320:26]
  assign _T_470 = ~ex_reg_ctrl_ren3 & ex_reg_inst[27]; // @[FPU.scala 784:53]
  assign _GEN_177 = {{1'd0}, _T_470}; // @[FPU.scala 784:36]
  assign _T_472 = ex_reg_ctrl_toint | ex_reg_ctrl_div; // @[FPU.scala 800:51]
  assign _T_473 = _T_472 | ex_reg_ctrl_sqrt; // @[FPU.scala 800:66]
  assign _T_474 = ex_reg_ctrl_fastpipe & ex_reg_ctrl_wflags; // @[FPU.scala 800:103]
  assign _T_475 = _T_473 | _T_474; // @[FPU.scala 800:82]
  assign _T_485 = {_T_383[22:0], 53'h0}; // @[FPU.scala 231:28]
  assign _GEN_178 = {{3'd0}, _T_383[31:23]}; // @[FPU.scala 234:31]
  assign _T_489 = _GEN_178 + 12'h800; // @[FPU.scala 234:31]
  assign _T_491 = _T_489 - 12'h100; // @[FPU.scala 234:48]
  assign _T_492 = _T_383[31:29] == 3'h0; // @[FPU.scala 235:19]
  assign _T_493 = _T_383[31:29] >= 3'h6; // @[FPU.scala 235:36]
  assign _T_494 = _T_492 | _T_493; // @[FPU.scala 235:25]
  assign _T_496 = {_T_383[31:29],_T_491[8:0]}; // @[Cat.scala 29:58]
  assign _T_498 = _T_494 ? _T_496 : _T_491; // @[FPU.scala 235:10]
  assign _T_500 = {_T_383[32],_T_498,_T_485[75:24]}; // @[Cat.scala 29:58]
  assign _T_505 = tag | _T_385; // @[package.scala 32:76]
  assign _T_507 = tag ? regfile_ex_rs_0_data : _T_500; // @[package.scala 32:76]
  assign _T_517 = {_T_412[22:0], 53'h0}; // @[FPU.scala 231:28]
  assign _GEN_179 = {{3'd0}, _T_412[31:23]}; // @[FPU.scala 234:31]
  assign _T_521 = _GEN_179 + 12'h800; // @[FPU.scala 234:31]
  assign _T_523 = _T_521 - 12'h100; // @[FPU.scala 234:48]
  assign _T_524 = _T_412[31:29] == 3'h0; // @[FPU.scala 235:19]
  assign _T_525 = _T_412[31:29] >= 3'h6; // @[FPU.scala 235:36]
  assign _T_526 = _T_524 | _T_525; // @[FPU.scala 235:25]
  assign _T_528 = {_T_412[31:29],_T_523[8:0]}; // @[Cat.scala 29:58]
  assign _T_530 = _T_526 ? _T_528 : _T_523; // @[FPU.scala 235:10]
  assign _T_532 = {_T_412[32],_T_530,_T_517[75:24]}; // @[Cat.scala 29:58]
  assign _T_537 = tag | _T_414; // @[package.scala 32:76]
  assign _T_539 = tag ? regfile_ex_rs_1_data : _T_532; // @[package.scala 32:76]
  assign _T_582 = {{1'd0}, io_fromint_data}; // @[FPU.scala 812:29]
  assign _T_682 = mem_ctrl_fma & mem_ctrl_singleOut; // @[FPU.scala 831:56]
  assign _T_683 = _T_682 ? 2'h2 : 2'h0; // @[FPU.scala 840:23]
  assign _T_685 = mem_ctrl_fma & ~mem_ctrl_singleOut; // @[FPU.scala 836:62]
  assign _T_686 = _T_685 ? 3'h4 : 3'h0; // @[FPU.scala 840:23]
  assign _T_687 = mem_ctrl_fastpipe | mem_ctrl_fromint; // @[FPU.scala 840:78]
  assign _GEN_186 = {{1'd0}, _T_687}; // @[FPU.scala 840:78]
  assign _T_688 = _GEN_186 | _T_683; // @[FPU.scala 840:78]
  assign _GEN_187 = {{1'd0}, _T_688}; // @[FPU.scala 840:78]
  assign memLatencyMask = _GEN_187 | _T_686; // @[FPU.scala 840:78]
  assign _T_689 = mem_ctrl_fma | mem_ctrl_fastpipe; // @[FPU.scala 856:48]
  assign _T_690 = _T_689 | mem_ctrl_fromint; // @[FPU.scala 856:69]
  assign mem_wen = mem_reg_valid & _T_690; // @[FPU.scala 856:31]
  assign _T_691 = ex_reg_ctrl_fastpipe ? 2'h2 : 2'h0; // @[FPU.scala 840:23]
  assign _T_692 = ex_reg_ctrl_fromint ? 2'h2 : 2'h0; // @[FPU.scala 840:23]
  assign _T_693 = ex_reg_ctrl_fma & ex_reg_ctrl_singleOut; // @[FPU.scala 831:56]
  assign _T_694 = _T_693 ? 3'h4 : 3'h0; // @[FPU.scala 840:23]
  assign _T_696 = ex_reg_ctrl_fma & ~ex_reg_ctrl_singleOut; // @[FPU.scala 836:62]
  assign _T_697 = _T_696 ? 4'h8 : 4'h0; // @[FPU.scala 840:23]
  assign _T_698 = _T_691 | _T_692; // @[FPU.scala 840:78]
  assign _GEN_188 = {{1'd0}, _T_698}; // @[FPU.scala 840:78]
  assign _T_699 = _GEN_188 | _T_694; // @[FPU.scala 840:78]
  assign _GEN_189 = {{1'd0}, _T_699}; // @[FPU.scala 840:78]
  assign _T_700 = _GEN_189 | _T_697; // @[FPU.scala 840:78]
  assign _GEN_190 = {{1'd0}, memLatencyMask}; // @[FPU.scala 857:62]
  assign _T_701 = _GEN_190 & _T_700; // @[FPU.scala 857:62]
  assign _T_702 = |_T_701; // @[FPU.scala 857:89]
  assign _T_703 = mem_wen & _T_702; // @[FPU.scala 857:43]
  assign _T_704 = ex_reg_ctrl_fastpipe ? 3'h4 : 3'h0; // @[FPU.scala 840:23]
  assign _T_705 = ex_reg_ctrl_fromint ? 3'h4 : 3'h0; // @[FPU.scala 840:23]
  assign _T_707 = _T_693 ? 4'h8 : 4'h0; // @[FPU.scala 840:23]
  assign _T_710 = _T_696 ? 5'h10 : 5'h0; // @[FPU.scala 840:23]
  assign _T_711 = _T_704 | _T_705; // @[FPU.scala 840:78]
  assign _GEN_191 = {{1'd0}, _T_711}; // @[FPU.scala 840:78]
  assign _T_712 = _GEN_191 | _T_707; // @[FPU.scala 840:78]
  assign _GEN_192 = {{1'd0}, _T_712}; // @[FPU.scala 840:78]
  assign _T_713 = _GEN_192 | _T_710; // @[FPU.scala 840:78]
  assign _GEN_193 = {{2'd0}, wen}; // @[FPU.scala 857:101]
  assign _T_714 = _GEN_193 & _T_713; // @[FPU.scala 857:101]
  assign _T_715 = |_T_714; // @[FPU.scala 857:128]
  assign _T_716 = _T_703 | _T_715; // @[FPU.scala 857:93]
  assign _GEN_194 = {{1'd0}, wen[2:1]}; // @[FPU.scala 866:23]
  assign _T_723 = _GEN_194 | memLatencyMask; // @[FPU.scala 866:23]
  assign _T_726 = ~write_port_busy & memLatencyMask[0]; // @[FPU.scala 869:30]
  assign _T_733 = _T_685 ? 2'h3 : 2'h0; // @[FPU.scala 842:63]
  assign _GEN_195 = {{1'd0}, mem_ctrl_fromint}; // @[FPU.scala 842:108]
  assign _T_735 = _GEN_195 | _T_683; // @[FPU.scala 842:108]
  assign _T_736 = _T_735 | _T_733; // @[FPU.scala 842:108]
  assign _T_740 = ~write_port_busy & memLatencyMask[1]; // @[FPU.scala 869:30]
  assign _T_754 = ~write_port_busy & memLatencyMask[2]; // @[FPU.scala 869:30]
  assign divSqrt_typeTag = divSqrt_1_io_outValid_div | divSqrt_1_io_outValid_sqrt; // @[FPU.scala 941:37]
  assign _T_1007 = divSqrt_io_outValid_div | divSqrt_io_outValid_sqrt; // @[FPU.scala 941:37]
  assign _GEN_156 = _T_1007 & ~divSqrt_killed; // @[FPU.scala 941:66]
  assign divSqrt_wen = divSqrt_typeTag ? ~divSqrt_killed : _GEN_156; // @[FPU.scala 941:66]
  assign wdouble = divSqrt_wen ? divSqrt_typeTag : ~wbInfo_0_single; // @[FPU.scala 879:20]
  assign _T_767 = wbInfo_0_pipeid == 2'h1; // @[package.scala 32:86]
  assign _T_768 = _T_767 ? ifpu_io_out_bits_data : fpmu_io_out_bits_data; // @[package.scala 32:76]
  assign _T_769 = wbInfo_0_pipeid == 2'h2; // @[package.scala 32:86]
  assign _T_770 = _T_769 ? sfma_io_out_bits_data : _T_768; // @[package.scala 32:76]
  assign _T_771 = wbInfo_0_pipeid == 2'h3; // @[package.scala 32:86]
  assign _T_772 = _T_771 ? dfma_io_out_bits_data : _T_770; // @[package.scala 32:76]
  assign _T_1023 = &divSqrt_1_io_out[63:61]; // @[FPU.scala 203:56]
  assign _T_1021 = divSqrt_1_io_out & 65'h1efefffffffffffff; // @[FPU.scala 361:25]
  assign _T_1024 = _T_1023 ? _T_1021 : divSqrt_1_io_out; // @[FPU.scala 362:10]
  assign _GEN_157 = divSqrt_io_out; // @[FPU.scala 941:66]
  assign divSqrt_wdata = divSqrt_typeTag ? _T_1024 : {{32'd0}, _GEN_157}; // @[FPU.scala 941:66]
  assign _T_773 = divSqrt_wen ? divSqrt_wdata : _T_772; // @[FPU.scala 880:22]
  assign _T_774 = &20'hfffff; // @[FPU.scala 286:42]
  assign _T_783 = {4'hf,_T_774,7'h7f,_T_773[31],20'hfffff,_T_773[32],_T_773[30:0]}; // @[Cat.scala 29:58]
  assign _T_784 = &3'h7; // @[FPU.scala 203:56]
  assign _T_785 = _T_784 ? _T_783 : 65'h1ffffffffffffffff; // @[FPU.scala 292:8]
  assign wdata_1 = wdouble ? _T_773 : _T_785; // @[package.scala 32:76]
  assign _T_789 = _T_767 ? ifpu_io_out_bits_exc : fpmu_io_out_bits_exc; // @[package.scala 32:76]
  assign _T_791 = _T_769 ? sfma_io_out_bits_exc : _T_789; // @[package.scala 32:76]
  assign wexc = _T_771 ? dfma_io_out_bits_exc : _T_791; // @[package.scala 32:76]
  assign frfWriteBundle_1_wrenf = wen[0] | divSqrt_wen; // @[FPU.scala 882:35]
  assign _T_807 = &wdata_1[63:61]; // @[FPU.scala 203:56]
  assign _T_811 = &wdata_1[51:32]; // @[FPU.scala 333:96]
  assign _T_812 = wdata_1[60] == _T_811; // @[FPU.scala 333:55]
  assign _T_813 = ~_T_807 | _T_812; // @[FPU.scala 333:31]
  assign _T_816 = _T_813 | reset; // @[FPU.scala 883:11]
  assign wb_toint_valid = wb_reg_valid & wb_ctrl_toint; // @[FPU.scala 898:37]
  assign _T_907 = wb_toint_valid | divSqrt_wen; // @[FPU.scala 900:41]
  assign _T_910 = wb_toint_valid ? wb_toint_exc : 5'h0; // @[FPU.scala 902:8]
  assign _GEN_158 = divSqrt_io_exceptionFlags; // @[FPU.scala 941:66]
  assign divSqrt_flags = divSqrt_typeTag ? divSqrt_1_io_exceptionFlags : _GEN_158; // @[FPU.scala 941:66]
  assign _T_911 = divSqrt_wen ? divSqrt_flags : 5'h0; // @[FPU.scala 903:8]
  assign _T_912 = _T_910 | _T_911; // @[FPU.scala 902:48]
  assign _T_914 = wen[0] ? wexc : 5'h0; // @[FPU.scala 904:8]
  assign _T_916 = mem_ctrl_div | mem_ctrl_sqrt; // @[FPU.scala 906:47]
  assign _T_917 = |wen; // @[FPU.scala 906:72]
  assign divSqrt_write_port_busy = _T_916 & _T_917; // @[FPU.scala 906:65]
  assign _T_918 = ex_reg_valid & ex_reg_ctrl_wflags; // @[FPU.scala 907:33]
  assign _T_919 = mem_reg_valid & mem_ctrl_wflags; // @[FPU.scala 907:68]
  assign _T_920 = _T_918 | _T_919; // @[FPU.scala 907:51]
  assign _T_922 = _T_920 | wb_toint_valid; // @[FPU.scala 907:87]
  assign _T_924 = _T_922 | _T_917; // @[FPU.scala 907:120]
  assign divSqrt_inFlight = ~divSqrt_1_io_inReady | ~divSqrt_io_inReady; // @[FPU.scala 934:34]
  assign _T_925 = _T_924 | divSqrt_inFlight; // @[FPU.scala 907:131]
  assign _T_927 = write_port_busy | divSqrt_write_port_busy; // @[FPU.scala 908:34]
  assign _T_934 = _T_685 | mem_ctrl_div; // @[FPU.scala 911:96]
  assign _T_942 = wen[0] & _T_771; // @[FPU.scala 912:60]
  assign _T_947 = io_inst[14:12] == 3'h5; // @[package.scala 15:47]
  assign _T_948 = io_inst[14:12] == 3'h6; // @[package.scala 15:47]
  assign _T_949 = _T_947 | _T_948; // @[package.scala 64:59]
  assign _T_951 = io_inst[14:12] == 3'h7; // @[FPU.scala 916:67]
  assign _T_952 = io_fcsr_rm >= 3'h5; // @[FPU.scala 916:87]
  assign _T_953 = _T_951 & _T_952; // @[FPU.scala 916:73]
  assign _T_961 = mem_reg_valid & mem_ctrl_singleOut; // @[FPU.scala 927:43]
  assign _T_963 = _T_961 & _T_916; // @[FPU.scala 927:65]
  assign _T_969 = {fpiu_io_out_bits_in_in1[51:0], 24'h0}; // @[FPU.scala 231:28]
  assign _T_973 = fpiu_io_out_bits_in_in1[63:52] + 12'h100; // @[FPU.scala 234:31]
  assign _T_975 = _T_973 - 12'h800; // @[FPU.scala 234:48]
  assign _T_976 = fpiu_io_out_bits_in_in1[63:61] == 3'h0; // @[FPU.scala 235:19]
  assign _T_977 = fpiu_io_out_bits_in_in1[63:61] >= 3'h6; // @[FPU.scala 235:36]
  assign _T_978 = _T_976 | _T_977; // @[FPU.scala 235:25]
  assign _T_980 = {fpiu_io_out_bits_in_in1[63:61],_T_975[5:0]}; // @[Cat.scala 29:58]
  assign _T_982 = _T_978 ? _T_980 : _T_975[8:0]; // @[FPU.scala 235:10]
  assign _T_983 = {fpiu_io_out_bits_in_in1[64],_T_982}; // @[Cat.scala 29:58]
  assign _T_988 = {fpiu_io_out_bits_in_in2[51:0], 24'h0}; // @[FPU.scala 231:28]
  assign _T_992 = fpiu_io_out_bits_in_in2[63:52] + 12'h100; // @[FPU.scala 234:31]
  assign _T_994 = _T_992 - 12'h800; // @[FPU.scala 234:48]
  assign _T_995 = fpiu_io_out_bits_in_in2[63:61] == 3'h0; // @[FPU.scala 235:19]
  assign _T_996 = fpiu_io_out_bits_in_in2[63:61] >= 3'h6; // @[FPU.scala 235:36]
  assign _T_997 = _T_995 | _T_996; // @[FPU.scala 235:25]
  assign _T_999 = {fpiu_io_out_bits_in_in2[63:61],_T_994[5:0]}; // @[Cat.scala 29:58]
  assign _T_1001 = _T_997 ? _T_999 : _T_994[8:0]; // @[FPU.scala 235:10]
  assign _T_1002 = {fpiu_io_out_bits_in_in2[64],_T_1001}; // @[Cat.scala 29:58]
  assign _T_1005 = divSqrt_io_inValid & divSqrt_io_inReady; // @[FPU.scala 936:32]
  assign _T_1010 = mem_reg_valid & ~mem_ctrl_singleOut; // @[FPU.scala 927:43]
  assign _T_1012 = _T_1010 & _T_916; // @[FPU.scala 927:65]
  assign _T_1016 = divSqrt_1_io_inValid & divSqrt_1_io_inReady; // @[FPU.scala 936:32]
  assign io_fcsr_flags_valid = _T_907 | wen[0]; // @[FPU.scala 900:23]
  assign io_fcsr_flags_bits = _T_912 | _T_914; // @[FPU.scala 901:22]
  assign io_store_data = fpiu_io_out_bits_store; // @[FPU.scala 802:17]
  assign io_toint_data = fpiu_io_out_bits_toint; // @[FPU.scala 803:17]
  assign io_fcsr_rdy = ~_T_925; // @[FPU.scala 907:15]
  assign io_nack_mem = _T_927 | divSqrt_inFlight; // @[FPU.scala 908:15]
  assign io_illegal_rm = _T_949 | _T_953; // @[FPU.scala 916:17]
  assign io_dec_wen = fp_decoder_io_sigs_wen; // @[FPU.scala 909:10]
  assign io_dec_ren1 = fp_decoder_io_sigs_ren1; // @[FPU.scala 909:10]
  assign io_dec_ren2 = fp_decoder_io_sigs_ren2; // @[FPU.scala 909:10]
  assign io_dec_ren3 = fp_decoder_io_sigs_ren3; // @[FPU.scala 909:10]
  assign io_sboard_set = wb_reg_valid & _T_936; // @[FPU.scala 911:17]
  assign io_sboard_clr = divSqrt_wen | _T_942; // @[FPU.scala 912:17]
  assign io_sboard_clra = divSqrt_wen ? divSqrt_waddr : wbInfo_0_rd; // @[FPU.scala 913:18]
  assign fp_decoder_io_inst = io_inst; // @[FPU.scala 695:22]
  assign sfma_clock = clock;
  assign sfma_reset = reset;
  assign sfma_io_in_valid = _T_377 & ex_reg_ctrl_singleOut; // @[FPU.scala 796:20]
  assign sfma_io_in_bits_ren3 = ex_reg_ctrl_ren3; // @[FPU.scala 797:19]
  assign sfma_io_in_bits_swap23 = ex_reg_ctrl_swap23; // @[FPU.scala 797:19]
  assign sfma_io_in_bits_rm = _T_375 ? io_fcsr_rm : ex_reg_inst[14:12]; // @[FPU.scala 797:19]
  assign sfma_io_in_bits_fmaCmd = ex_reg_inst[3:2] | _GEN_177; // @[FPU.scala 797:19]
  assign sfma_io_in_bits_in1 = {{32'd0}, _T_407}; // @[FPU.scala 797:19]
  assign sfma_io_in_bits_in2 = {{32'd0}, _T_436}; // @[FPU.scala 797:19]
  assign sfma_io_in_bits_in3 = {{32'd0}, _T_465}; // @[FPU.scala 797:19]
  assign fpiu_clock = clock;
  assign fpiu_io_in_valid = ex_reg_valid & _T_475; // @[FPU.scala 800:20]
  assign fpiu_io_in_bits_ren2 = ex_reg_ctrl_ren2; // @[FPU.scala 801:19]
  assign fpiu_io_in_bits_singleIn = ex_reg_ctrl_singleIn; // @[FPU.scala 801:19]
  assign fpiu_io_in_bits_singleOut = ex_reg_ctrl_singleOut; // @[FPU.scala 801:19]
  assign fpiu_io_in_bits_wflags = ex_reg_ctrl_wflags; // @[FPU.scala 801:19]
  assign fpiu_io_in_bits_rm = _T_375 ? io_fcsr_rm : ex_reg_inst[14:12]; // @[FPU.scala 801:19]
  assign fpiu_io_in_bits_typ = ex_reg_inst[21:20]; // @[FPU.scala 801:19]
  assign fpiu_io_in_bits_in1 = _T_505 ? _T_507 : 65'he008000000000000; // @[FPU.scala 801:19]
  assign fpiu_io_in_bits_in2 = _T_537 ? _T_539 : 65'he008000000000000; // @[FPU.scala 801:19]
  assign ifpu_clock = clock;
  assign ifpu_reset = reset;
  assign ifpu_io_in_valid = ex_reg_valid & ex_reg_ctrl_fromint; // @[FPU.scala 810:20]
  assign ifpu_io_in_bits_singleIn = fpiu_io_in_bits_singleIn; // @[FPU.scala 811:19]
  assign ifpu_io_in_bits_wflags = fpiu_io_in_bits_wflags; // @[FPU.scala 811:19]
  assign ifpu_io_in_bits_rm = fpiu_io_in_bits_rm; // @[FPU.scala 811:19]
  assign ifpu_io_in_bits_typ = fpiu_io_in_bits_typ; // @[FPU.scala 811:19]
  assign ifpu_io_in_bits_in1 = _T_582[63:0]; // @[FPU.scala 811:19 FPU.scala 812:23]
  assign fpmu_clock = clock;
  assign fpmu_reset = reset;
  assign fpmu_io_in_valid = ex_reg_valid & ex_reg_ctrl_fastpipe; // @[FPU.scala 815:20]
  assign fpmu_io_in_bits_ren2 = fpiu_io_in_bits_ren2; // @[FPU.scala 816:19]
  assign fpmu_io_in_bits_singleOut = fpiu_io_in_bits_singleOut; // @[FPU.scala 816:19]
  assign fpmu_io_in_bits_wflags = fpiu_io_in_bits_wflags; // @[FPU.scala 816:19]
  assign fpmu_io_in_bits_rm = fpiu_io_in_bits_rm; // @[FPU.scala 816:19]
  assign fpmu_io_in_bits_in1 = fpiu_io_in_bits_in1; // @[FPU.scala 816:19]
  assign fpmu_io_in_bits_in2 = fpiu_io_in_bits_in2; // @[FPU.scala 816:19]
  assign fpmu_io_lt = fpiu_io_out_bits_lt; // @[FPU.scala 817:14]
  assign dfma_clock = clock;
  assign dfma_reset = reset;
  assign dfma_io_in_valid = _T_377 & ~ex_reg_ctrl_singleOut; // @[FPU.scala 834:28]
  assign dfma_io_in_bits_ren3 = ex_reg_ctrl_ren3; // @[FPU.scala 835:27]
  assign dfma_io_in_bits_swap23 = ex_reg_ctrl_swap23; // @[FPU.scala 835:27]
  assign dfma_io_in_bits_rm = _T_375 ? io_fcsr_rm : ex_reg_inst[14:12]; // @[FPU.scala 835:27]
  assign dfma_io_in_bits_fmaCmd = ex_reg_inst[3:2] | _GEN_177; // @[FPU.scala 835:27]
  assign dfma_io_in_bits_in1 = regfile_ex_rs_0_data; // @[FPU.scala 835:27]
  assign dfma_io_in_bits_in2 = regfile_ex_rs_1_data; // @[FPU.scala 835:27]
  assign dfma_io_in_bits_in3 = regfile_ex_rs_2_data; // @[FPU.scala 835:27]
  assign divSqrt_clock = clock;
  assign divSqrt_reset = reset;
  assign divSqrt_io_inValid = _T_963 & ~divSqrt_inFlight; // @[FPU.scala 927:26]
  assign divSqrt_io_sqrtOp = mem_ctrl_sqrt; // @[FPU.scala 928:25]
  assign divSqrt_io_a = {_T_983,_T_969[75:53]}; // @[FPU.scala 929:20]
  assign divSqrt_io_b = {_T_1002,_T_988[75:53]}; // @[FPU.scala 930:20]
  assign divSqrt_io_roundingMode = fpiu_io_out_bits_in_rm; // @[FPU.scala 931:31]
  assign divSqrt_1_clock = clock;
  assign divSqrt_1_reset = reset;
  assign divSqrt_1_io_inValid = _T_1012 & ~divSqrt_inFlight; // @[FPU.scala 927:26]
  assign divSqrt_1_io_sqrtOp = mem_ctrl_sqrt; // @[FPU.scala 928:25]
  assign divSqrt_1_io_a = fpiu_io_out_bits_in_in1; // @[FPU.scala 929:20]
  assign divSqrt_1_io_b = fpiu_io_out_bits_in_in2; // @[FPU.scala 930:20]
  assign divSqrt_1_io_roundingMode = fpiu_io_out_bits_in_rm; // @[FPU.scala 931:31]
  assign FPU_cov_read_addr = FPU_state;
  assign FPU_cov_read_data = FPU_cov[FPU_cov_read_addr]; // @[Coverage map for FPU]
  assign FPU_cov_write_data = 1'h1;
  assign FPU_cov_write_addr = FPU_state;
  assign FPU_cov_write_mask = 1'h1;
  assign FPU_cov_write_en = 1'h1;
  assign wbInfo_0_single_shl = wbInfo_0_single;
  assign wbInfo_0_single_pad = {19'h0,wbInfo_0_single_shl};
  assign ex_reg_ctrl_fromint_shl = {ex_reg_ctrl_fromint, 16'h0};
  assign ex_reg_ctrl_fromint_pad = {3'h0,ex_reg_ctrl_fromint_shl};
  assign wb_ctrl_toint_shl = {wb_ctrl_toint, 19'h0};
  assign wb_ctrl_toint_pad = wb_ctrl_toint_shl;
  assign ex_reg_ctrl_fastpipe_shl = {ex_reg_ctrl_fastpipe, 13'h0};
  assign ex_reg_ctrl_fastpipe_pad = {6'h0,ex_reg_ctrl_fastpipe_shl};
  assign mem_reg_valid_shl = {mem_reg_valid, 1'h0};
  assign mem_reg_valid_pad = {18'h0,mem_reg_valid_shl};
  assign write_port_busy_shl = {write_port_busy, 14'h0};
  assign write_port_busy_pad = {5'h0,write_port_busy_shl};
  assign ex_reg_ctrl_singleIn_shl = {ex_reg_ctrl_singleIn, 2'h0};
  assign ex_reg_ctrl_singleIn_pad = {17'h0,ex_reg_ctrl_singleIn_shl};
  assign mem_ctrl_fastpipe_shl = {mem_ctrl_fastpipe, 1'h0};
  assign mem_ctrl_fastpipe_pad = {18'h0,mem_ctrl_fastpipe_shl};
  assign wbInfo_0_pipeid_shl = {wbInfo_0_pipeid, 12'h0};
  assign wbInfo_0_pipeid_pad = {6'h0,wbInfo_0_pipeid_shl};
  assign load_wb_double_shl = {load_wb_double, 1'h0};
  assign load_wb_double_pad = {18'h0,load_wb_double_shl};
  assign ex_reg_ctrl_singleOut_shl = ex_reg_ctrl_singleOut;
  assign ex_reg_ctrl_singleOut_pad = {19'h0,ex_reg_ctrl_singleOut_shl};
  assign wen_shl = {wen, 1'h0};
  assign wen_pad = {16'h0,wen_shl};
  assign mem_ctrl_toint_shl = {mem_ctrl_toint, 14'h0};
  assign mem_ctrl_toint_pad = {5'h0,mem_ctrl_toint_shl};
  assign wb_reg_valid_shl = {wb_reg_valid, 7'h0};
  assign wb_reg_valid_pad = {12'h0,wb_reg_valid_shl};
  assign ex_reg_ctrl_fma_shl = {ex_reg_ctrl_fma, 2'h0};
  assign ex_reg_ctrl_fma_pad = {17'h0,ex_reg_ctrl_fma_shl};
  assign mem_ctrl_singleOut_shl = {mem_ctrl_singleOut, 4'h0};
  assign mem_ctrl_singleOut_pad = {15'h0,mem_ctrl_singleOut_shl};
  assign mem_ctrl_fromint_shl = {mem_ctrl_fromint, 8'h0};
  assign mem_ctrl_fromint_pad = {11'h0,mem_ctrl_fromint_shl};
  assign mem_ctrl_fma_shl = {mem_ctrl_fma, 17'h0};
  assign mem_ctrl_fma_pad = {2'h0,mem_ctrl_fma_shl};
  assign ex_reg_valid_shl = {ex_reg_valid, 7'h0};
  assign ex_reg_valid_pad = {12'h0,ex_reg_valid_shl};
  assign divSqrt_killed_shl = {divSqrt_killed, 16'h0};
  assign divSqrt_killed_pad = {3'h0,divSqrt_killed_shl};
  assign FPU_xor7 = wbInfo_0_single_pad ^ ex_reg_ctrl_fromint_pad;
  assign FPU_xor18 = ex_reg_ctrl_fastpipe_pad ^ mem_reg_valid_pad;
  assign FPU_xor8 = wb_ctrl_toint_pad ^ FPU_xor18;
  assign FPU_xor3 = FPU_xor7 ^ FPU_xor8;
  assign FPU_xor9 = write_port_busy_pad ^ ex_reg_ctrl_singleIn_pad;
  assign FPU_xor22 = wbInfo_0_pipeid_pad ^ load_wb_double_pad;
  assign FPU_xor10 = mem_ctrl_fastpipe_pad ^ FPU_xor22;
  assign FPU_xor4 = FPU_xor9 ^ FPU_xor10;
  assign FPU_xor1 = FPU_xor3 ^ FPU_xor4;
  assign FPU_xor11 = ex_reg_ctrl_singleOut_pad ^ wen_pad;
  assign FPU_xor26 = wb_reg_valid_pad ^ ex_reg_ctrl_fma_pad;
  assign FPU_xor12 = mem_ctrl_toint_pad ^ FPU_xor26;
  assign FPU_xor5 = FPU_xor11 ^ FPU_xor12;
  assign FPU_xor13 = mem_ctrl_singleOut_pad ^ mem_ctrl_fromint_pad;
  assign FPU_xor30 = ex_reg_valid_pad ^ divSqrt_killed_pad;
  assign FPU_xor14 = mem_ctrl_fma_pad ^ FPU_xor30;
  assign FPU_xor6 = FPU_xor13 ^ FPU_xor14;
  assign FPU_xor2 = FPU_xor5 ^ FPU_xor6;
  assign FPU_xor0 = FPU_xor1 ^ FPU_xor2;
  assign divSqrt_1_sum = FPU_covSum + divSqrt_1_io_covSum;
  assign ifpu_sum = divSqrt_1_sum + ifpu_io_covSum;
  assign divSqrt_sum = ifpu_sum + divSqrt_io_covSum;
  assign fpmu_sum = divSqrt_sum + fpmu_io_covSum;
  assign fp_decoder_sum = fpmu_sum + fp_decoder_io_covSum;
  assign dfma_sum = fp_decoder_sum + dfma_io_covSum;
  assign fpiu_sum = dfma_sum + fpiu_io_covSum;
  assign sfma_sum = fpiu_sum + sfma_io_covSum;
  assign io_covSum = sfma_sum;
  assign stopEn0 = load_wb & ~_T_271;
  assign stopEn1 = frfWriteBundle_1_wrenf & ~_T_816;
  assign divSqrt_metaAssert_wire = divSqrt_metaAssert;
  assign dfma_metaAssert_wire = dfma_metaAssert;
  assign fpiu_metaAssert_wire = fpiu_metaAssert;
  assign fpmu_metaAssert_wire = fpmu_metaAssert;
  assign divSqrt_1_metaAssert_wire = divSqrt_1_metaAssert;
  assign sfma_metaAssert_wire = sfma_metaAssert;
  assign ifpu_metaAssert_wire = ifpu_metaAssert;
  assign fp_decoder_metaAssert_wire = fp_decoder_metaAssert;
  assign FPU_or3 = stopEn0 | stopEn1;
  assign FPU_or10 = divSqrt_metaAssert_wire | divSqrt_1_metaAssert_wire;
  assign FPU_or4 = fp_decoder_metaAssert_wire | FPU_or10;
  assign FPU_or1 = FPU_or3 | FPU_or4;
  assign FPU_or5 = fpiu_metaAssert_wire | dfma_metaAssert_wire;
  assign FPU_or14 = ifpu_metaAssert_wire | sfma_metaAssert_wire;
  assign FPU_or6 = fpmu_metaAssert_wire | FPU_or14;
  assign FPU_or2 = FPU_or5 | FPU_or6;
  assign FPU_or0 = FPU_or1 | FPU_or2;
  assign metaAssert = FPU_metaAssert;
  assign divSqrt_1_metaReset = metaReset | divSqrt_1_halt;
  assign ifpu_metaReset = metaReset | ifpu_halt;
  assign divSqrt_metaReset = metaReset | divSqrt_halt;
  assign fpmu_metaReset = metaReset | fpmu_halt;
  assign dfma_metaReset = metaReset | dfma_halt;
  assign fpiu_metaReset = metaReset | fpiu_halt;
  assign sfma_metaReset = metaReset | sfma_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {3{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regfile[initvar] = _RAND_0[64:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ex_reg_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ex_reg_inst = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ex_reg_ctrl_ren2 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ex_reg_ctrl_ren3 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ex_reg_ctrl_swap23 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ex_reg_ctrl_singleIn = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ex_reg_ctrl_singleOut = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ex_reg_ctrl_fromint = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  ex_reg_ctrl_toint = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  ex_reg_ctrl_fastpipe = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  ex_reg_ctrl_fma = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  ex_reg_ctrl_div = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  ex_reg_ctrl_sqrt = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  ex_reg_ctrl_wflags = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  ex_ra_0 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  ex_ra_1 = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  ex_ra_2 = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  load_wb = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  load_wb_double = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  load_wb_data = _RAND_20[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  load_wb_tag = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mem_reg_valid = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mem_reg_inst = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  wb_reg_valid = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  mem_ctrl_singleOut = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mem_ctrl_fromint = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mem_ctrl_toint = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  mem_ctrl_fastpipe = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  mem_ctrl_fma = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  mem_ctrl_div = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  mem_ctrl_sqrt = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  mem_ctrl_wflags = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  wb_ctrl_toint = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  divSqrt_waddr = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  wen = _RAND_35[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  wbInfo_0_rd = _RAND_36[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  wbInfo_0_single = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  wbInfo_0_pipeid = _RAND_38[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  wbInfo_1_rd = _RAND_39[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  wbInfo_1_single = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  wbInfo_1_pipeid = _RAND_41[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  wbInfo_2_rd = _RAND_42[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  wbInfo_2_single = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  wbInfo_2_pipeid = _RAND_44[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  write_port_busy = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  divSqrt_killed = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  wb_toint_exc = _RAND_47[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_936 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  FPU_state = _RAND_49[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    FPU_cov[initvar] = _RAND_50[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  FPU_covSum = _RAND_51[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  FPU_metaAssert = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(regfile__T_251_en & regfile__T_251_mask) begin
      regfile[regfile__T_251_addr] <= regfile__T_251_data; // @[FPU.scala 748:20]
    end
    if(regfile__T_818_en & regfile__T_818_mask) begin
      regfile[regfile__T_818_addr] <= regfile__T_818_data; // @[FPU.scala 748:20]
    end
    if (metaReset) begin
      ex_reg_valid <= 1'h0;
    end else if (reset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= io_valid;
    end
    if (metaReset) begin
      ex_reg_inst <= 32'h0;
    end else if (io_valid) begin
      ex_reg_inst <= io_inst;
    end
    if (metaReset) begin
      ex_reg_ctrl_ren2 <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_ren2 <= fp_decoder_io_sigs_ren2;
    end
    if (metaReset) begin
      ex_reg_ctrl_ren3 <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_ren3 <= fp_decoder_io_sigs_ren3;
    end
    if (metaReset) begin
      ex_reg_ctrl_swap23 <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_swap23 <= fp_decoder_io_sigs_swap23;
    end
    if (metaReset) begin
      ex_reg_ctrl_singleIn <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_singleIn <= fp_decoder_io_sigs_singleIn;
    end
    if (metaReset) begin
      ex_reg_ctrl_singleOut <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_singleOut <= fp_decoder_io_sigs_singleOut;
    end
    if (metaReset) begin
      ex_reg_ctrl_fromint <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_fromint <= fp_decoder_io_sigs_fromint;
    end
    if (metaReset) begin
      ex_reg_ctrl_toint <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_toint <= fp_decoder_io_sigs_toint;
    end
    if (metaReset) begin
      ex_reg_ctrl_fastpipe <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_fastpipe <= fp_decoder_io_sigs_fastpipe;
    end
    if (metaReset) begin
      ex_reg_ctrl_fma <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_fma <= fp_decoder_io_sigs_fma;
    end
    if (metaReset) begin
      ex_reg_ctrl_div <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_div <= fp_decoder_io_sigs_div;
    end
    if (metaReset) begin
      ex_reg_ctrl_sqrt <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_sqrt <= fp_decoder_io_sigs_sqrt;
    end
    if (metaReset) begin
      ex_reg_ctrl_wflags <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_wflags <= fp_decoder_io_sigs_wflags;
    end
    if (metaReset) begin
      ex_ra_0 <= 5'h0;
    end else if (io_valid) begin
      if (fp_decoder_io_sigs_ren2) begin
        if (fp_decoder_io_sigs_swap12) begin
          ex_ra_0 <= io_inst[24:20];
        end else if (fp_decoder_io_sigs_ren1) begin
          if (~fp_decoder_io_sigs_swap12) begin
            ex_ra_0 <= io_inst[19:15];
          end
        end
      end else if (fp_decoder_io_sigs_ren1) begin
        if (~fp_decoder_io_sigs_swap12) begin
          ex_ra_0 <= io_inst[19:15];
        end
      end
    end
    if (metaReset) begin
      ex_ra_1 <= 5'h0;
    end else if (io_valid) begin
      if (fp_decoder_io_sigs_ren2) begin
        if (_T_371) begin
          ex_ra_1 <= io_inst[24:20];
        end else if (fp_decoder_io_sigs_ren1) begin
          if (fp_decoder_io_sigs_swap12) begin
            ex_ra_1 <= io_inst[19:15];
          end
        end
      end else if (fp_decoder_io_sigs_ren1) begin
        if (fp_decoder_io_sigs_swap12) begin
          ex_ra_1 <= io_inst[19:15];
        end
      end
    end
    if (metaReset) begin
      ex_ra_2 <= 5'h0;
    end else if (io_valid) begin
      if (fp_decoder_io_sigs_ren3) begin
        ex_ra_2 <= io_inst[31:27];
      end else if (fp_decoder_io_sigs_ren2) begin
        if (fp_decoder_io_sigs_swap23) begin
          ex_ra_2 <= io_inst[24:20];
        end
      end
    end
    if (metaReset) begin
      load_wb <= 1'h0;
    end else begin
      load_wb <= io_dmem_resp_val;
    end
    if (metaReset) begin
      load_wb_double <= 1'h0;
    end else if (io_dmem_resp_val) begin
      load_wb_double <= io_dmem_resp_type[0];
    end
    if (metaReset) begin
      load_wb_data <= 64'h0;
    end else if (io_dmem_resp_val) begin
      load_wb_data <= io_dmem_resp_data;
    end
    if (metaReset) begin
      load_wb_tag <= 5'h0;
    end else if (io_dmem_resp_val) begin
      load_wb_tag <= io_dmem_resp_tag;
    end
    if (metaReset) begin
      mem_reg_valid <= 1'h0;
    end else if (reset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= _T_5;
    end
    if (metaReset) begin
      mem_reg_inst <= 32'h0;
    end else if (ex_reg_valid) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if (metaReset) begin
      wb_reg_valid <= 1'h0;
    end else if (reset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= _T_9;
    end
    if (metaReset) begin
      mem_ctrl_singleOut <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_singleOut <= ex_reg_ctrl_singleOut;
    end
    if (metaReset) begin
      mem_ctrl_fromint <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_fromint <= ex_reg_ctrl_fromint;
    end
    if (metaReset) begin
      mem_ctrl_toint <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_toint <= ex_reg_ctrl_toint;
    end
    if (metaReset) begin
      mem_ctrl_fastpipe <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_fastpipe <= ex_reg_ctrl_fastpipe;
    end
    if (metaReset) begin
      mem_ctrl_fma <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_fma <= ex_reg_ctrl_fma;
    end
    if (metaReset) begin
      mem_ctrl_div <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_div <= ex_reg_ctrl_div;
    end
    if (metaReset) begin
      mem_ctrl_sqrt <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_sqrt <= ex_reg_ctrl_sqrt;
    end
    if (metaReset) begin
      mem_ctrl_wflags <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_wflags <= ex_reg_ctrl_wflags;
    end
    if (metaReset) begin
      wb_ctrl_toint <= 1'h0;
    end else if (mem_reg_valid) begin
      wb_ctrl_toint <= mem_ctrl_toint;
    end
    if (metaReset) begin
      divSqrt_waddr <= 5'h0;
    end else if (_T_1016) begin
      divSqrt_waddr <= mem_reg_inst[11:7];
    end else if (_T_1005) begin
      divSqrt_waddr <= mem_reg_inst[11:7];
    end
    if (metaReset) begin
      wen <= 3'h0;
    end else if (reset) begin
      wen <= 3'h0;
    end else if (mem_wen) begin
      if (~killm) begin
        wen <= _T_723;
      end else begin
        wen <= {{1'd0}, wen[2:1]};
      end
    end else begin
      wen <= {{1'd0}, wen[2:1]};
    end
    if (metaReset) begin
      wbInfo_0_rd <= 5'h0;
    end else if (mem_wen) begin
      if (_T_726) begin
        wbInfo_0_rd <= mem_reg_inst[11:7];
      end else if (wen[1]) begin
        wbInfo_0_rd <= wbInfo_1_rd;
      end
    end else if (wen[1]) begin
      wbInfo_0_rd <= wbInfo_1_rd;
    end
    if (metaReset) begin
      wbInfo_0_single <= 1'h0;
    end else if (mem_wen) begin
      if (_T_726) begin
        wbInfo_0_single <= mem_ctrl_singleOut;
      end else if (wen[1]) begin
        wbInfo_0_single <= wbInfo_1_single;
      end
    end else if (wen[1]) begin
      wbInfo_0_single <= wbInfo_1_single;
    end
    if (metaReset) begin
      wbInfo_0_pipeid <= 2'h0;
    end else if (mem_wen) begin
      if (_T_726) begin
        wbInfo_0_pipeid <= _T_736;
      end else if (wen[1]) begin
        wbInfo_0_pipeid <= wbInfo_1_pipeid;
      end
    end else if (wen[1]) begin
      wbInfo_0_pipeid <= wbInfo_1_pipeid;
    end
    if (metaReset) begin
      wbInfo_1_rd <= 5'h0;
    end else if (mem_wen) begin
      if (_T_740) begin
        wbInfo_1_rd <= mem_reg_inst[11:7];
      end else if (wen[2]) begin
        wbInfo_1_rd <= wbInfo_2_rd;
      end
    end else if (wen[2]) begin
      wbInfo_1_rd <= wbInfo_2_rd;
    end
    if (metaReset) begin
      wbInfo_1_single <= 1'h0;
    end else if (mem_wen) begin
      if (_T_740) begin
        wbInfo_1_single <= mem_ctrl_singleOut;
      end else if (wen[2]) begin
        wbInfo_1_single <= wbInfo_2_single;
      end
    end else if (wen[2]) begin
      wbInfo_1_single <= wbInfo_2_single;
    end
    if (metaReset) begin
      wbInfo_1_pipeid <= 2'h0;
    end else if (mem_wen) begin
      if (_T_740) begin
        wbInfo_1_pipeid <= _T_736;
      end else if (wen[2]) begin
        wbInfo_1_pipeid <= wbInfo_2_pipeid;
      end
    end else if (wen[2]) begin
      wbInfo_1_pipeid <= wbInfo_2_pipeid;
    end
    if (metaReset) begin
      wbInfo_2_rd <= 5'h0;
    end else if (mem_wen) begin
      if (_T_754) begin
        wbInfo_2_rd <= mem_reg_inst[11:7];
      end
    end
    if (metaReset) begin
      wbInfo_2_single <= 1'h0;
    end else if (mem_wen) begin
      if (_T_754) begin
        wbInfo_2_single <= mem_ctrl_singleOut;
      end
    end
    if (metaReset) begin
      wbInfo_2_pipeid <= 2'h0;
    end else if (mem_wen) begin
      if (_T_754) begin
        wbInfo_2_pipeid <= _T_736;
      end
    end
    if (metaReset) begin
      write_port_busy <= 1'h0;
    end else if (ex_reg_valid) begin
      write_port_busy <= _T_716;
    end
    if (metaReset) begin
      divSqrt_killed <= 1'h0;
    end else if (_T_1016) begin
      divSqrt_killed <= killm;
    end else if (_T_1005) begin
      divSqrt_killed <= killm;
    end
    if (metaReset) begin
      wb_toint_exc <= 5'h0;
    end else if (mem_ctrl_toint) begin
      wb_toint_exc <= fpiu_io_out_bits_exc;
    end
    if (metaReset) begin
      _T_936 <= 1'h0;
    end else begin
      _T_936 <= _T_934 | mem_ctrl_sqrt;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (load_wb & ~_T_271) begin
          $fwrite(32'h80000002,"Assertion failed\n    at FPU.scala:752 assert(consistent(wdata))\n"); // @[FPU.scala 752:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (load_wb & ~_T_271) begin
          $fatal; // @[FPU.scala 752:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (frfWriteBundle_1_wrenf & ~_T_816) begin
          $fwrite(32'h80000002,"Assertion failed\n    at FPU.scala:883 assert(consistent(wdata))\n"); // @[FPU.scala 883:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (frfWriteBundle_1_wrenf & ~_T_816) begin
          $fatal; // @[FPU.scala 883:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    FPU_state <= FPU_xor0;
    if (!(FPU_cov_read_data)) begin
      FPU_covSum <= FPU_covSum + 1'h1;
    end
    if (metaReset) begin
      FPU_metaAssert <= 1'h0;
    end else begin
      FPU_metaAssert <= FPU_metaAssert | FPU_or0;
    end
  end
  always @(posedge clock) begin
    if(FPU_cov_write_en & FPU_cov_write_mask) begin
      FPU_cov[FPU_cov_write_addr] <= FPU_cov_write_data; // @[Coverage map for FPU]
    end
  end
endmodule
module HellaCacheArbiter(
  input         clock,
  output        io_requestor_0_req_ready,
  input         io_requestor_0_req_valid,
  input  [39:0] io_requestor_0_req_bits_addr,
  input         io_requestor_0_s1_kill,
  output        io_requestor_0_s2_nack,
  output        io_requestor_0_resp_valid,
  output [63:0] io_requestor_0_resp_bits_data,
  output        io_requestor_0_s2_xcpt_ae_ld,
  output        io_requestor_1_req_ready,
  input         io_requestor_1_req_valid,
  input  [39:0] io_requestor_1_req_bits_addr,
  input  [6:0]  io_requestor_1_req_bits_tag,
  input  [4:0]  io_requestor_1_req_bits_cmd,
  input  [1:0]  io_requestor_1_req_bits_size,
  input         io_requestor_1_req_bits_signed,
  input         io_requestor_1_s1_kill,
  input  [63:0] io_requestor_1_s1_data_data,
  output        io_requestor_1_s2_nack,
  output        io_requestor_1_resp_valid,
  output [6:0]  io_requestor_1_resp_bits_tag,
  output [1:0]  io_requestor_1_resp_bits_size,
  output [63:0] io_requestor_1_resp_bits_data,
  output        io_requestor_1_resp_bits_replay,
  output        io_requestor_1_resp_bits_has_data,
  output [63:0] io_requestor_1_resp_bits_data_word_bypass,
  output        io_requestor_1_replay_next,
  output        io_requestor_1_s2_xcpt_ma_ld,
  output        io_requestor_1_s2_xcpt_ma_st,
  output        io_requestor_1_s2_xcpt_pf_ld,
  output        io_requestor_1_s2_xcpt_pf_st,
  output        io_requestor_1_s2_xcpt_ae_ld,
  output        io_requestor_1_s2_xcpt_ae_st,
  output        io_requestor_1_ordered,
  output        io_requestor_1_perf_release,
  output        io_requestor_1_perf_grant,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output [6:0]  io_mem_req_bits_tag,
  output [4:0]  io_mem_req_bits_cmd,
  output [1:0]  io_mem_req_bits_size,
  output        io_mem_req_bits_signed,
  output        io_mem_req_bits_phys,
  output        io_mem_s1_kill,
  output [63:0] io_mem_s1_data_data,
  input         io_mem_s2_nack,
  input         io_mem_resp_valid,
  input  [6:0]  io_mem_resp_bits_tag,
  input  [1:0]  io_mem_resp_bits_size,
  input  [63:0] io_mem_resp_bits_data,
  input         io_mem_resp_bits_replay,
  input         io_mem_resp_bits_has_data,
  input  [63:0] io_mem_resp_bits_data_word_bypass,
  input         io_mem_replay_next,
  input         io_mem_s2_xcpt_ma_ld,
  input         io_mem_s2_xcpt_ma_st,
  input         io_mem_s2_xcpt_pf_ld,
  input         io_mem_s2_xcpt_pf_st,
  input         io_mem_s2_xcpt_ae_ld,
  input         io_mem_s2_xcpt_ae_st,
  input         io_mem_ordered,
  input         io_mem_perf_release,
  input         io_mem_perf_grant,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  _T; // @[HellaCacheArbiter.scala 19:20]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[HellaCacheArbiter.scala 20:20]
  reg [31:0] _RAND_1;
  wire [7:0] _T_6; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1; // @[HellaCacheArbiter.scala 49:26]
  reg  HellaCacheArbiter_state; // @[Register tracking HellaCacheArbiter state]
  reg [31:0] _RAND_2;
  reg  HellaCacheArbiter_cov [0:1]; // @[Coverage map for HellaCacheArbiter]
  reg [31:0] _RAND_3;
  wire  HellaCacheArbiter_cov_read_data; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_read_addr; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_write_data; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_write_addr; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_write_mask; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_write_en; // @[Coverage map for HellaCacheArbiter]
  reg [29:0] HellaCacheArbiter_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_4;
  wire  _T_shl;
  wire  _T_pad;
  assign _T_6 = {io_requestor_1_req_bits_tag,1'h1}; // @[Cat.scala 29:58]
  assign _GEN_1 = io_requestor_0_req_valid ? 8'h0 : _T_6; // @[HellaCacheArbiter.scala 49:26]
  assign io_requestor_0_req_ready = io_mem_req_ready; // @[HellaCacheArbiter.scala 25:31]
  assign io_requestor_0_s2_nack = io_mem_s2_nack & ~_T_1; // @[HellaCacheArbiter.scala 64:31]
  assign io_requestor_0_resp_valid = io_mem_resp_valid & ~io_mem_resp_bits_tag[0]; // @[HellaCacheArbiter.scala 60:18]
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data; // @[HellaCacheArbiter.scala 69:17]
  assign io_requestor_0_s2_xcpt_ae_ld = io_mem_s2_xcpt_ae_ld; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_req_ready = io_requestor_0_req_ready & ~io_requestor_0_req_valid; // @[HellaCacheArbiter.scala 27:33]
  assign io_requestor_1_s2_nack = io_mem_s2_nack & _T_1; // @[HellaCacheArbiter.scala 64:31]
  assign io_requestor_1_resp_valid = io_mem_resp_valid & io_mem_resp_bits_tag[0]; // @[HellaCacheArbiter.scala 60:18]
  assign io_requestor_1_resp_bits_tag = {{1'd0}, io_mem_resp_bits_tag[6:1]}; // @[HellaCacheArbiter.scala 69:17 HellaCacheArbiter.scala 70:21]
  assign io_requestor_1_resp_bits_size = io_mem_resp_bits_size; // @[HellaCacheArbiter.scala 69:17]
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data; // @[HellaCacheArbiter.scala 69:17]
  assign io_requestor_1_resp_bits_replay = io_mem_resp_bits_replay; // @[HellaCacheArbiter.scala 69:17]
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data; // @[HellaCacheArbiter.scala 69:17]
  assign io_requestor_1_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass; // @[HellaCacheArbiter.scala 69:17]
  assign io_requestor_1_replay_next = io_mem_replay_next; // @[HellaCacheArbiter.scala 72:35]
  assign io_requestor_1_s2_xcpt_ma_ld = io_mem_s2_xcpt_ma_ld; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_s2_xcpt_ma_st = io_mem_s2_xcpt_ma_st; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_s2_xcpt_pf_ld = io_mem_s2_xcpt_pf_ld; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_s2_xcpt_pf_st = io_mem_s2_xcpt_pf_st; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_s2_xcpt_ae_ld = io_mem_s2_xcpt_ae_ld; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_s2_xcpt_ae_st = io_mem_s2_xcpt_ae_st; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_ordered = io_mem_ordered; // @[HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_perf_release = io_mem_perf_release; // @[HellaCacheArbiter.scala 63:28]
  assign io_requestor_1_perf_grant = io_mem_perf_grant; // @[HellaCacheArbiter.scala 63:28]
  assign io_mem_req_valid = io_requestor_0_req_valid | io_requestor_1_req_valid; // @[HellaCacheArbiter.scala 24:22]
  assign io_mem_req_bits_addr = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr; // @[HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 32:25]
  assign io_mem_req_bits_tag = _GEN_1[6:0]; // @[HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 33:29 HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 33:29]
  assign io_mem_req_bits_cmd = io_requestor_0_req_valid ? 5'h0 : io_requestor_1_req_bits_cmd; // @[HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 32:25]
  assign io_mem_req_bits_size = io_requestor_0_req_valid ? 2'h3 : io_requestor_1_req_bits_size; // @[HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 32:25]
  assign io_mem_req_bits_signed = io_requestor_0_req_valid ? 1'h0 : io_requestor_1_req_bits_signed; // @[HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 32:25]
  assign io_mem_req_bits_phys = io_requestor_0_req_valid; // @[HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 32:25]
  assign io_mem_s1_kill = _T ? io_requestor_1_s1_kill : io_requestor_0_s1_kill; // @[HellaCacheArbiter.scala 37:24 HellaCacheArbiter.scala 37:24]
  assign io_mem_s1_data_data = _T ? io_requestor_1_s1_data_data : 64'h0; // @[HellaCacheArbiter.scala 38:24 HellaCacheArbiter.scala 38:24]
  assign HellaCacheArbiter_cov_read_addr = HellaCacheArbiter_state;
  assign HellaCacheArbiter_cov_read_data = HellaCacheArbiter_cov[HellaCacheArbiter_cov_read_addr]; // @[Coverage map for HellaCacheArbiter]
  assign HellaCacheArbiter_cov_write_data = 1'h1;
  assign HellaCacheArbiter_cov_write_addr = HellaCacheArbiter_state;
  assign HellaCacheArbiter_cov_write_mask = 1'h1;
  assign HellaCacheArbiter_cov_write_en = 1'h1;
  assign _T_shl = _T;
  assign _T_pad = _T_shl;
  assign io_covSum = HellaCacheArbiter_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  HellaCacheArbiter_state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    HellaCacheArbiter_cov[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  HellaCacheArbiter_covSum = _RAND_4[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T <= 1'h0;
    end else if (io_requestor_0_req_valid) begin
      _T <= 1'h0;
    end else begin
      _T <= 1'h1;
    end
    if (metaReset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= _T;
    end
    HellaCacheArbiter_state <= _T_pad;
    if (!(HellaCacheArbiter_cov_read_data)) begin
      HellaCacheArbiter_covSum <= HellaCacheArbiter_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(HellaCacheArbiter_cov_write_en & HellaCacheArbiter_cov_write_mask) begin
      HellaCacheArbiter_cov[HellaCacheArbiter_cov_write_addr] <= HellaCacheArbiter_cov_write_data; // @[Coverage map for HellaCacheArbiter]
    end
  end
endmodule
module PTW(
  input         clock,
  input         reset,
  output        io_requestor_0_req_ready,
  input         io_requestor_0_req_valid,
  input  [26:0] io_requestor_0_req_bits_bits_addr,
  output        io_requestor_0_resp_valid,
  output        io_requestor_0_resp_bits_ae,
  output [53:0] io_requestor_0_resp_bits_pte_ppn,
  output        io_requestor_0_resp_bits_pte_d,
  output        io_requestor_0_resp_bits_pte_a,
  output        io_requestor_0_resp_bits_pte_g,
  output        io_requestor_0_resp_bits_pte_u,
  output        io_requestor_0_resp_bits_pte_x,
  output        io_requestor_0_resp_bits_pte_w,
  output        io_requestor_0_resp_bits_pte_r,
  output        io_requestor_0_resp_bits_pte_v,
  output [1:0]  io_requestor_0_resp_bits_level,
  output        io_requestor_0_resp_bits_homogeneous,
  output [3:0]  io_requestor_0_ptbr_mode,
  output        io_requestor_0_status_debug,
  output [1:0]  io_requestor_0_status_dprv,
  output        io_requestor_0_status_mxr,
  output        io_requestor_0_status_sum,
  output        io_requestor_0_pmp_0_cfg_l,
  output [1:0]  io_requestor_0_pmp_0_cfg_a,
  output        io_requestor_0_pmp_0_cfg_x,
  output        io_requestor_0_pmp_0_cfg_w,
  output        io_requestor_0_pmp_0_cfg_r,
  output [29:0] io_requestor_0_pmp_0_addr,
  output [31:0] io_requestor_0_pmp_0_mask,
  output        io_requestor_0_pmp_1_cfg_l,
  output [1:0]  io_requestor_0_pmp_1_cfg_a,
  output        io_requestor_0_pmp_1_cfg_x,
  output        io_requestor_0_pmp_1_cfg_w,
  output        io_requestor_0_pmp_1_cfg_r,
  output [29:0] io_requestor_0_pmp_1_addr,
  output [31:0] io_requestor_0_pmp_1_mask,
  output        io_requestor_0_pmp_2_cfg_l,
  output [1:0]  io_requestor_0_pmp_2_cfg_a,
  output        io_requestor_0_pmp_2_cfg_x,
  output        io_requestor_0_pmp_2_cfg_w,
  output        io_requestor_0_pmp_2_cfg_r,
  output [29:0] io_requestor_0_pmp_2_addr,
  output [31:0] io_requestor_0_pmp_2_mask,
  output        io_requestor_0_pmp_3_cfg_l,
  output [1:0]  io_requestor_0_pmp_3_cfg_a,
  output        io_requestor_0_pmp_3_cfg_x,
  output        io_requestor_0_pmp_3_cfg_w,
  output        io_requestor_0_pmp_3_cfg_r,
  output [29:0] io_requestor_0_pmp_3_addr,
  output [31:0] io_requestor_0_pmp_3_mask,
  output        io_requestor_0_pmp_4_cfg_l,
  output [1:0]  io_requestor_0_pmp_4_cfg_a,
  output        io_requestor_0_pmp_4_cfg_x,
  output        io_requestor_0_pmp_4_cfg_w,
  output        io_requestor_0_pmp_4_cfg_r,
  output [29:0] io_requestor_0_pmp_4_addr,
  output [31:0] io_requestor_0_pmp_4_mask,
  output        io_requestor_0_pmp_5_cfg_l,
  output [1:0]  io_requestor_0_pmp_5_cfg_a,
  output        io_requestor_0_pmp_5_cfg_x,
  output        io_requestor_0_pmp_5_cfg_w,
  output        io_requestor_0_pmp_5_cfg_r,
  output [29:0] io_requestor_0_pmp_5_addr,
  output [31:0] io_requestor_0_pmp_5_mask,
  output        io_requestor_0_pmp_6_cfg_l,
  output [1:0]  io_requestor_0_pmp_6_cfg_a,
  output        io_requestor_0_pmp_6_cfg_x,
  output        io_requestor_0_pmp_6_cfg_w,
  output        io_requestor_0_pmp_6_cfg_r,
  output [29:0] io_requestor_0_pmp_6_addr,
  output [31:0] io_requestor_0_pmp_6_mask,
  output        io_requestor_0_pmp_7_cfg_l,
  output [1:0]  io_requestor_0_pmp_7_cfg_a,
  output        io_requestor_0_pmp_7_cfg_x,
  output        io_requestor_0_pmp_7_cfg_w,
  output        io_requestor_0_pmp_7_cfg_r,
  output [29:0] io_requestor_0_pmp_7_addr,
  output [31:0] io_requestor_0_pmp_7_mask,
  output        io_requestor_1_req_ready,
  input         io_requestor_1_req_valid,
  input         io_requestor_1_req_bits_valid,
  input  [26:0] io_requestor_1_req_bits_bits_addr,
  output        io_requestor_1_resp_valid,
  output        io_requestor_1_resp_bits_ae,
  output [53:0] io_requestor_1_resp_bits_pte_ppn,
  output        io_requestor_1_resp_bits_pte_d,
  output        io_requestor_1_resp_bits_pte_a,
  output        io_requestor_1_resp_bits_pte_g,
  output        io_requestor_1_resp_bits_pte_u,
  output        io_requestor_1_resp_bits_pte_x,
  output        io_requestor_1_resp_bits_pte_w,
  output        io_requestor_1_resp_bits_pte_r,
  output        io_requestor_1_resp_bits_pte_v,
  output [1:0]  io_requestor_1_resp_bits_level,
  output        io_requestor_1_resp_bits_homogeneous,
  output [3:0]  io_requestor_1_ptbr_mode,
  output        io_requestor_1_status_debug,
  output [1:0]  io_requestor_1_status_prv,
  output        io_requestor_1_pmp_0_cfg_l,
  output [1:0]  io_requestor_1_pmp_0_cfg_a,
  output        io_requestor_1_pmp_0_cfg_x,
  output        io_requestor_1_pmp_0_cfg_w,
  output        io_requestor_1_pmp_0_cfg_r,
  output [29:0] io_requestor_1_pmp_0_addr,
  output [31:0] io_requestor_1_pmp_0_mask,
  output        io_requestor_1_pmp_1_cfg_l,
  output [1:0]  io_requestor_1_pmp_1_cfg_a,
  output        io_requestor_1_pmp_1_cfg_x,
  output        io_requestor_1_pmp_1_cfg_w,
  output        io_requestor_1_pmp_1_cfg_r,
  output [29:0] io_requestor_1_pmp_1_addr,
  output [31:0] io_requestor_1_pmp_1_mask,
  output        io_requestor_1_pmp_2_cfg_l,
  output [1:0]  io_requestor_1_pmp_2_cfg_a,
  output        io_requestor_1_pmp_2_cfg_x,
  output        io_requestor_1_pmp_2_cfg_w,
  output        io_requestor_1_pmp_2_cfg_r,
  output [29:0] io_requestor_1_pmp_2_addr,
  output [31:0] io_requestor_1_pmp_2_mask,
  output        io_requestor_1_pmp_3_cfg_l,
  output [1:0]  io_requestor_1_pmp_3_cfg_a,
  output        io_requestor_1_pmp_3_cfg_x,
  output        io_requestor_1_pmp_3_cfg_w,
  output        io_requestor_1_pmp_3_cfg_r,
  output [29:0] io_requestor_1_pmp_3_addr,
  output [31:0] io_requestor_1_pmp_3_mask,
  output        io_requestor_1_pmp_4_cfg_l,
  output [1:0]  io_requestor_1_pmp_4_cfg_a,
  output        io_requestor_1_pmp_4_cfg_x,
  output        io_requestor_1_pmp_4_cfg_w,
  output        io_requestor_1_pmp_4_cfg_r,
  output [29:0] io_requestor_1_pmp_4_addr,
  output [31:0] io_requestor_1_pmp_4_mask,
  output        io_requestor_1_pmp_5_cfg_l,
  output [1:0]  io_requestor_1_pmp_5_cfg_a,
  output        io_requestor_1_pmp_5_cfg_x,
  output        io_requestor_1_pmp_5_cfg_w,
  output        io_requestor_1_pmp_5_cfg_r,
  output [29:0] io_requestor_1_pmp_5_addr,
  output [31:0] io_requestor_1_pmp_5_mask,
  output        io_requestor_1_pmp_6_cfg_l,
  output [1:0]  io_requestor_1_pmp_6_cfg_a,
  output        io_requestor_1_pmp_6_cfg_x,
  output        io_requestor_1_pmp_6_cfg_w,
  output        io_requestor_1_pmp_6_cfg_r,
  output [29:0] io_requestor_1_pmp_6_addr,
  output [31:0] io_requestor_1_pmp_6_mask,
  output        io_requestor_1_pmp_7_cfg_l,
  output [1:0]  io_requestor_1_pmp_7_cfg_a,
  output        io_requestor_1_pmp_7_cfg_x,
  output        io_requestor_1_pmp_7_cfg_w,
  output        io_requestor_1_pmp_7_cfg_r,
  output [29:0] io_requestor_1_pmp_7_addr,
  output [31:0] io_requestor_1_pmp_7_mask,
  output [63:0] io_requestor_1_customCSRs_csrs_0_value,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output        io_mem_s1_kill,
  input         io_mem_s2_nack,
  input         io_mem_resp_valid,
  input  [63:0] io_mem_resp_bits_data,
  input         io_mem_s2_xcpt_ae_ld,
  input  [3:0]  io_dpath_ptbr_mode,
  input  [43:0] io_dpath_ptbr_ppn,
  input         io_dpath_sfence_valid,
  input         io_dpath_sfence_bits_rs1,
  input         io_dpath_status_debug,
  input  [1:0]  io_dpath_status_dprv,
  input  [1:0]  io_dpath_status_prv,
  input         io_dpath_status_mxr,
  input         io_dpath_status_sum,
  input         io_dpath_pmp_0_cfg_l,
  input  [1:0]  io_dpath_pmp_0_cfg_a,
  input         io_dpath_pmp_0_cfg_x,
  input         io_dpath_pmp_0_cfg_w,
  input         io_dpath_pmp_0_cfg_r,
  input  [29:0] io_dpath_pmp_0_addr,
  input  [31:0] io_dpath_pmp_0_mask,
  input         io_dpath_pmp_1_cfg_l,
  input  [1:0]  io_dpath_pmp_1_cfg_a,
  input         io_dpath_pmp_1_cfg_x,
  input         io_dpath_pmp_1_cfg_w,
  input         io_dpath_pmp_1_cfg_r,
  input  [29:0] io_dpath_pmp_1_addr,
  input  [31:0] io_dpath_pmp_1_mask,
  input         io_dpath_pmp_2_cfg_l,
  input  [1:0]  io_dpath_pmp_2_cfg_a,
  input         io_dpath_pmp_2_cfg_x,
  input         io_dpath_pmp_2_cfg_w,
  input         io_dpath_pmp_2_cfg_r,
  input  [29:0] io_dpath_pmp_2_addr,
  input  [31:0] io_dpath_pmp_2_mask,
  input         io_dpath_pmp_3_cfg_l,
  input  [1:0]  io_dpath_pmp_3_cfg_a,
  input         io_dpath_pmp_3_cfg_x,
  input         io_dpath_pmp_3_cfg_w,
  input         io_dpath_pmp_3_cfg_r,
  input  [29:0] io_dpath_pmp_3_addr,
  input  [31:0] io_dpath_pmp_3_mask,
  input         io_dpath_pmp_4_cfg_l,
  input  [1:0]  io_dpath_pmp_4_cfg_a,
  input         io_dpath_pmp_4_cfg_x,
  input         io_dpath_pmp_4_cfg_w,
  input         io_dpath_pmp_4_cfg_r,
  input  [29:0] io_dpath_pmp_4_addr,
  input  [31:0] io_dpath_pmp_4_mask,
  input         io_dpath_pmp_5_cfg_l,
  input  [1:0]  io_dpath_pmp_5_cfg_a,
  input         io_dpath_pmp_5_cfg_x,
  input         io_dpath_pmp_5_cfg_w,
  input         io_dpath_pmp_5_cfg_r,
  input  [29:0] io_dpath_pmp_5_addr,
  input  [31:0] io_dpath_pmp_5_mask,
  input         io_dpath_pmp_6_cfg_l,
  input  [1:0]  io_dpath_pmp_6_cfg_a,
  input         io_dpath_pmp_6_cfg_x,
  input         io_dpath_pmp_6_cfg_w,
  input         io_dpath_pmp_6_cfg_r,
  input  [29:0] io_dpath_pmp_6_addr,
  input  [31:0] io_dpath_pmp_6_mask,
  input         io_dpath_pmp_7_cfg_l,
  input  [1:0]  io_dpath_pmp_7_cfg_a,
  input         io_dpath_pmp_7_cfg_x,
  input         io_dpath_pmp_7_cfg_w,
  input         io_dpath_pmp_7_cfg_r,
  input  [29:0] io_dpath_pmp_7_addr,
  input  [31:0] io_dpath_pmp_7_mask,
  input  [63:0] io_dpath_customCSRs_csrs_0_value,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  output [19:0] Checking_PTW_regstate,			//Jaewon_PTW_regstate
  output [29:0] Checking_PTW_covSum				//Jaewon_PTW_regstate
  );
  assign Checking_PTW_regstate = PTW_state; 	//Jaewon_PTW_regstate
  assign Checking_PTW_covSum = PTW_covSum; 		//Jaewon_PTW_regstate
  wire  arb_io_in_0_ready; // @[PTW.scala 105:19]
  wire  arb_io_in_0_valid; // @[PTW.scala 105:19]
  wire [26:0] arb_io_in_0_bits_bits_addr; // @[PTW.scala 105:19]
  wire  arb_io_in_1_ready; // @[PTW.scala 105:19]
  wire  arb_io_in_1_valid; // @[PTW.scala 105:19]
  wire  arb_io_in_1_bits_valid; // @[PTW.scala 105:19]
  wire [26:0] arb_io_in_1_bits_bits_addr; // @[PTW.scala 105:19]
  wire  arb_io_out_ready; // @[PTW.scala 105:19]
  wire  arb_io_out_valid; // @[PTW.scala 105:19]
  wire  arb_io_out_bits_valid; // @[PTW.scala 105:19]
  wire [26:0] arb_io_out_bits_bits_addr; // @[PTW.scala 105:19]
  wire  arb_io_chosen; // @[PTW.scala 105:19]
  wire [29:0] arb_io_covSum; // @[PTW.scala 105:19]
  wire  arb_metaAssert; // @[PTW.scala 105:19]
  wire [2:0] OptimizationBarrier_io_x; // @[package.scala 236:25]
  wire [2:0] OptimizationBarrier_io_y; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_metaAssert; // @[package.scala 236:25]
  wire [53:0] OptimizationBarrier_1_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_d; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_a; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_g; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_x; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_w; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_r; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_v; // @[package.scala 236:25]
  wire [53:0] OptimizationBarrier_1_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_d; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_a; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_g; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_x; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_w; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_r; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_v; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_1_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_metaAssert; // @[package.scala 236:25]
  reg [2:0] state; // @[PTW.scala 103:18]
  reg [31:0] _RAND_0;
  reg  resp_valid_0; // @[PTW.scala 109:23]
  reg [31:0] _RAND_1;
  reg  resp_valid_1; // @[PTW.scala 109:23]
  reg [31:0] _RAND_2;
  wire  _T_2; // @[PTW.scala 111:24]
  reg  invalidated; // @[PTW.scala 118:24]
  reg [31:0] _RAND_3;
  reg [1:0] count; // @[PTW.scala 119:18]
  reg [31:0] _RAND_4;
  reg  resp_ae; // @[PTW.scala 120:24]
  reg [31:0] _RAND_5;
  reg [26:0] r_req_addr; // @[PTW.scala 123:18]
  reg [31:0] _RAND_6;
  reg  r_req_dest; // @[PTW.scala 124:23]
  reg [31:0] _RAND_7;
  reg [53:0] r_pte_ppn; // @[PTW.scala 125:18]
  reg [63:0] _RAND_8;
  reg  r_pte_d; // @[PTW.scala 125:18]
  reg [31:0] _RAND_9;
  reg  r_pte_a; // @[PTW.scala 125:18]
  reg [31:0] _RAND_10;
  reg  r_pte_g; // @[PTW.scala 125:18]
  reg [31:0] _RAND_11;
  reg  r_pte_u; // @[PTW.scala 125:18]
  reg [31:0] _RAND_12;
  reg  r_pte_x; // @[PTW.scala 125:18]
  reg [31:0] _RAND_13;
  reg  r_pte_w; // @[PTW.scala 125:18]
  reg [31:0] _RAND_14;
  reg  r_pte_r; // @[PTW.scala 125:18]
  reg [31:0] _RAND_15;
  reg  r_pte_v; // @[PTW.scala 125:18]
  reg [31:0] _RAND_16;
  reg  mem_resp_valid; // @[PTW.scala 127:31]
  reg [31:0] _RAND_17;
  reg [63:0] mem_resp_data; // @[PTW.scala 128:30]
  reg [63:0] _RAND_18;
  wire  tmp_v; // @[PTW.scala 139:33]
  wire  tmp_r; // @[PTW.scala 139:33]
  wire  tmp_w; // @[PTW.scala 139:33]
  wire  tmp_x; // @[PTW.scala 139:33]
  wire  tmp_u; // @[PTW.scala 139:33]
  wire  tmp_g; // @[PTW.scala 139:33]
  wire  tmp_a; // @[PTW.scala 139:33]
  wire  tmp_d; // @[PTW.scala 139:33]
  wire [53:0] tmp_ppn; // @[PTW.scala 139:33]
  wire  _T_19; // @[PTW.scala 142:17]
  wire  _T_20; // @[PTW.scala 142:26]
  wire  _T_21; // @[PTW.scala 145:21]
  wire  _T_23; // @[PTW.scala 145:95]
  wire  _T_24; // @[PTW.scala 145:26]
  wire  _GEN_0; // @[PTW.scala 145:102]
  wire  _T_25; // @[PTW.scala 145:21]
  wire  _T_27; // @[PTW.scala 145:95]
  wire  _T_28; // @[PTW.scala 145:26]
  wire  _GEN_1; // @[PTW.scala 145:102]
  wire  res_v; // @[PTW.scala 142:36]
  wire  invalid_paddr; // @[PTW.scala 147:32]
  wire  _T_31; // @[PTW.scala 68:33]
  wire  _T_33; // @[PTW.scala 68:39]
  wire  _T_35; // @[PTW.scala 68:45]
  wire  _T_37; // @[PTW.scala 149:30]
  wire  _T_38; // @[PTW.scala 149:57]
  wire  traverse; // @[PTW.scala 149:48]
  wire [8:0] vpn_idxs_0; // @[PTW.scala 151:60]
  wire [8:0] vpn_idxs_1; // @[PTW.scala 151:90]
  wire [8:0] vpn_idxs_2; // @[PTW.scala 151:90]
  wire  _T_42; // @[package.scala 32:86]
  wire [8:0] _T_43; // @[package.scala 32:76]
  wire  _T_44; // @[package.scala 32:86]
  wire [8:0] _T_45; // @[package.scala 32:76]
  wire  _T_46; // @[package.scala 32:86]
  wire [8:0] vpn_idx; // @[package.scala 32:76]
  wire [62:0] _T_47; // @[Cat.scala 29:58]
  wire [65:0] pte_addr; // @[PTW.scala 153:29]
  wire [53:0] choices_0; // @[Cat.scala 29:58]
  wire [53:0] choices_1; // @[Cat.scala 29:58]
  wire [53:0] fragmented_superpage_ppn; // @[package.scala 32:76]
  wire  _T_55; // @[Decoupled.scala 40:37]
  reg [6:0] _T_56; // @[Replacement.scala 158:30]
  reg [31:0] _RAND_19;
  reg [7:0] valid; // @[PTW.scala 168:24]
  reg [31:0] _RAND_20;
  reg [31:0] tags_0; // @[PTW.scala 169:19]
  reg [31:0] _RAND_21;
  reg [31:0] tags_1; // @[PTW.scala 169:19]
  reg [31:0] _RAND_22;
  reg [31:0] tags_2; // @[PTW.scala 169:19]
  reg [31:0] _RAND_23;
  reg [31:0] tags_3; // @[PTW.scala 169:19]
  reg [31:0] _RAND_24;
  reg [31:0] tags_4; // @[PTW.scala 169:19]
  reg [31:0] _RAND_25;
  reg [31:0] tags_5; // @[PTW.scala 169:19]
  reg [31:0] _RAND_26;
  reg [31:0] tags_6; // @[PTW.scala 169:19]
  reg [31:0] _RAND_27;
  reg [31:0] tags_7; // @[PTW.scala 169:19]
  reg [31:0] _RAND_28;
  reg [19:0] data_0; // @[PTW.scala 170:19]
  reg [31:0] _RAND_29;
  reg [19:0] data_1; // @[PTW.scala 170:19]
  reg [31:0] _RAND_30;
  reg [19:0] data_2; // @[PTW.scala 170:19]
  reg [31:0] _RAND_31;
  reg [19:0] data_3; // @[PTW.scala 170:19]
  reg [31:0] _RAND_32;
  reg [19:0] data_4; // @[PTW.scala 170:19]
  reg [31:0] _RAND_33;
  reg [19:0] data_5; // @[PTW.scala 170:19]
  reg [31:0] _RAND_34;
  reg [19:0] data_6; // @[PTW.scala 170:19]
  reg [31:0] _RAND_35;
  reg [19:0] data_7; // @[PTW.scala 170:19]
  reg [31:0] _RAND_36;
  wire [65:0] _GEN_108; // @[PTW.scala 172:27]
  wire  _T_57; // @[PTW.scala 172:27]
  wire [65:0] _GEN_109; // @[PTW.scala 172:27]
  wire  _T_58; // @[PTW.scala 172:27]
  wire [65:0] _GEN_110; // @[PTW.scala 172:27]
  wire  _T_59; // @[PTW.scala 172:27]
  wire [65:0] _GEN_111; // @[PTW.scala 172:27]
  wire  _T_60; // @[PTW.scala 172:27]
  wire [65:0] _GEN_112; // @[PTW.scala 172:27]
  wire  _T_61; // @[PTW.scala 172:27]
  wire [65:0] _GEN_113; // @[PTW.scala 172:27]
  wire  _T_62; // @[PTW.scala 172:27]
  wire [65:0] _GEN_114; // @[PTW.scala 172:27]
  wire  _T_63; // @[PTW.scala 172:27]
  wire [65:0] _GEN_115; // @[PTW.scala 172:27]
  wire  _T_64; // @[PTW.scala 172:27]
  wire [7:0] _T_71; // @[Cat.scala 29:58]
  wire [7:0] hits; // @[PTW.scala 172:48]
  wire  hit; // @[PTW.scala 173:20]
  wire  _T_72; // @[PTW.scala 174:26]
  wire  _T_74; // @[PTW.scala 174:38]
  wire  _T_76; // @[PTW.scala 174:46]
  wire  _T_77; // @[PTW.scala 175:25]
  wire  _T_86; // @[Replacement.scala 240:16]
  wire [1:0] _T_87; // @[Cat.scala 29:58]
  wire  _T_93; // @[Replacement.scala 240:16]
  wire [1:0] _T_94; // @[Cat.scala 29:58]
  wire [1:0] _T_95; // @[Replacement.scala 240:16]
  wire [2:0] _T_96; // @[Cat.scala 29:58]
  wire  _T_98; // @[OneHot.scala 47:40]
  wire  _T_99; // @[OneHot.scala 47:40]
  wire  _T_100; // @[OneHot.scala 47:40]
  wire  _T_101; // @[OneHot.scala 47:40]
  wire  _T_102; // @[OneHot.scala 47:40]
  wire  _T_103; // @[OneHot.scala 47:40]
  wire  _T_104; // @[OneHot.scala 47:40]
  wire [2:0] _T_106; // @[Mux.scala 47:69]
  wire [2:0] _T_107; // @[Mux.scala 47:69]
  wire [2:0] _T_108; // @[Mux.scala 47:69]
  wire [2:0] _T_109; // @[Mux.scala 47:69]
  wire [2:0] _T_110; // @[Mux.scala 47:69]
  wire [2:0] _T_111; // @[Mux.scala 47:69]
  wire [2:0] _T_112; // @[Mux.scala 47:69]
  wire [2:0] r; // @[PTW.scala 175:18]
  wire [7:0] _T_113; // @[OneHot.scala 58:35]
  wire [7:0] _T_114; // @[PTW.scala 176:22]
  wire [53:0] res_ppn; // @[PTW.scala 141:13]
  wire  _T_115; // @[PTW.scala 180:24]
  wire  _T_116; // @[PTW.scala 180:15]
  wire  _T_119; // @[OneHot.scala 32:14]
  wire [3:0] _T_120; // @[OneHot.scala 32:28]
  wire  _T_123; // @[OneHot.scala 32:14]
  wire [1:0] _T_124; // @[OneHot.scala 32:28]
  wire [2:0] _T_127; // @[Cat.scala 29:58]
  wire  _T_141; // @[Replacement.scala 193:16]
  wire  _T_145; // @[Replacement.scala 196:16]
  wire [2:0] _T_147; // @[Cat.scala 29:58]
  wire [2:0] _T_148; // @[Replacement.scala 193:16]
  wire  _T_157; // @[Replacement.scala 193:16]
  wire  _T_161; // @[Replacement.scala 196:16]
  wire [2:0] _T_163; // @[Cat.scala 29:58]
  wire [2:0] _T_164; // @[Replacement.scala 196:16]
  wire [6:0] _T_166; // @[Cat.scala 29:58]
  wire  _T_168; // @[PTW.scala 181:33]
  wire  pte_cache_hit; // @[PTW.scala 186:10]
  wire [19:0] _T_186; // @[Mux.scala 27:72]
  wire [19:0] _T_187; // @[Mux.scala 27:72]
  wire [19:0] _T_188; // @[Mux.scala 27:72]
  wire [19:0] _T_189; // @[Mux.scala 27:72]
  wire [19:0] _T_190; // @[Mux.scala 27:72]
  wire [19:0] _T_191; // @[Mux.scala 27:72]
  wire [19:0] _T_192; // @[Mux.scala 27:72]
  wire [19:0] _T_193; // @[Mux.scala 27:72]
  wire [19:0] _T_194; // @[Mux.scala 27:72]
  wire [19:0] _T_195; // @[Mux.scala 27:72]
  wire [19:0] _T_196; // @[Mux.scala 27:72]
  wire [19:0] _T_197; // @[Mux.scala 27:72]
  wire [19:0] _T_198; // @[Mux.scala 27:72]
  wire [19:0] _T_199; // @[Mux.scala 27:72]
  wire [19:0] pte_cache_data; // @[Mux.scala 27:72]
  wire  _T_202; // @[PTW.scala 245:56]
  wire  _T_205; // @[PTW.scala 247:48]
  wire [65:0] _T_215; // @[Parameters.scala 137:31]
  wire [66:0] _T_216; // @[Parameters.scala 137:49]
  wire [66:0] _T_218; // @[Parameters.scala 137:52]
  wire  _T_219; // @[Parameters.scala 137:67]
  wire [65:0] _T_220; // @[Parameters.scala 137:31]
  wire [66:0] _T_221; // @[Parameters.scala 137:49]
  wire [66:0] _T_223; // @[Parameters.scala 137:52]
  wire  _T_224; // @[Parameters.scala 137:67]
  wire [65:0] _T_225; // @[Parameters.scala 137:31]
  wire [66:0] _T_226; // @[Parameters.scala 137:49]
  wire [66:0] _T_228; // @[Parameters.scala 137:52]
  wire  _T_229; // @[Parameters.scala 137:67]
  wire  _T_231; // @[TLBPermissions.scala 98:65]
  wire  pmaPgLevelHomogeneous_1; // @[TLBPermissions.scala 98:65]
  wire [66:0] _T_235; // @[Parameters.scala 137:49]
  wire [66:0] _T_262; // @[Parameters.scala 137:52]
  wire  _T_263; // @[Parameters.scala 137:67]
  wire [65:0] _T_264; // @[Parameters.scala 137:31]
  wire [66:0] _T_265; // @[Parameters.scala 137:49]
  wire [66:0] _T_267; // @[Parameters.scala 137:52]
  wire  _T_268; // @[Parameters.scala 137:67]
  wire [65:0] _T_269; // @[Parameters.scala 137:31]
  wire [66:0] _T_270; // @[Parameters.scala 137:49]
  wire [66:0] _T_272; // @[Parameters.scala 137:52]
  wire  _T_273; // @[Parameters.scala 137:67]
  wire [65:0] _T_274; // @[Parameters.scala 137:31]
  wire [66:0] _T_275; // @[Parameters.scala 137:49]
  wire [66:0] _T_277; // @[Parameters.scala 137:52]
  wire  _T_278; // @[Parameters.scala 137:67]
  wire  _T_295; // @[TLBPermissions.scala 98:65]
  wire  _T_296; // @[TLBPermissions.scala 98:65]
  wire  _T_297; // @[TLBPermissions.scala 98:65]
  wire  _T_298; // @[TLBPermissions.scala 98:65]
  wire  _T_299; // @[TLBPermissions.scala 98:65]
  wire  pmaPgLevelHomogeneous_2; // @[TLBPermissions.scala 98:65]
  wire  _T_352; // @[package.scala 32:76]
  wire  _T_354; // @[package.scala 32:76]
  wire  pmaHomogeneous; // @[package.scala 32:76]
  wire [65:0] _T_357; // @[PTW.scala 268:92]
  wire  _T_364; // @[package.scala 32:76]
  wire  _T_366; // @[package.scala 32:76]
  wire  _T_368; // @[package.scala 32:76]
  wire [31:0] _T_369; // @[PMP.scala 62:36]
  wire [31:0] _T_371; // @[PMP.scala 62:48]
  wire [65:0] _GEN_116; // @[PMP.scala 100:53]
  wire [65:0] _T_373; // @[PMP.scala 100:53]
  wire  _T_375; // @[PMP.scala 100:78]
  wire  _T_382; // @[PMP.scala 100:78]
  wire  _T_389; // @[PMP.scala 100:78]
  wire  _T_391; // @[package.scala 32:76]
  wire  _T_393; // @[package.scala 32:76]
  wire  _T_395; // @[package.scala 32:76]
  wire  _T_396; // @[PMP.scala 100:21]
  wire  _T_409; // @[PMP.scala 109:32]
  wire [31:0] _T_412; // @[package.scala 32:76]
  wire [31:0] _T_414; // @[package.scala 32:76]
  wire [31:0] _T_416; // @[package.scala 32:76]
  wire [65:0] _GEN_120; // @[PMP.scala 112:30]
  wire [65:0] _T_417; // @[PMP.scala 112:30]
  wire [31:0] _T_429; // @[PMP.scala 113:53]
  wire [65:0] _GEN_122; // @[PMP.scala 113:40]
  wire  _T_430; // @[PMP.scala 113:40]
  wire  _T_433; // @[PMP.scala 115:41]
  wire  _T_434; // @[PMP.scala 120:58]
  wire  _T_435; // @[PMP.scala 120:8]
  wire  _T_442; // @[package.scala 32:76]
  wire  _T_444; // @[package.scala 32:76]
  wire  _T_446; // @[package.scala 32:76]
  wire [31:0] _T_447; // @[PMP.scala 62:36]
  wire [31:0] _T_449; // @[PMP.scala 62:48]
  wire [65:0] _GEN_123; // @[PMP.scala 100:53]
  wire [65:0] _T_451; // @[PMP.scala 100:53]
  wire  _T_453; // @[PMP.scala 100:78]
  wire  _T_460; // @[PMP.scala 100:78]
  wire  _T_467; // @[PMP.scala 100:78]
  wire  _T_469; // @[package.scala 32:76]
  wire  _T_471; // @[package.scala 32:76]
  wire  _T_473; // @[package.scala 32:76]
  wire  _T_474; // @[PMP.scala 100:21]
  wire  _T_487; // @[PMP.scala 109:32]
  wire [31:0] _T_507; // @[PMP.scala 113:53]
  wire [65:0] _GEN_131; // @[PMP.scala 113:40]
  wire  _T_508; // @[PMP.scala 113:40]
  wire  _T_509; // @[PMP.scala 115:21]
  wire  _T_510; // @[PMP.scala 115:62]
  wire  _T_511; // @[PMP.scala 115:41]
  wire  _T_512; // @[PMP.scala 120:58]
  wire  _T_513; // @[PMP.scala 120:8]
  wire  _T_514; // @[PMP.scala 140:10]
  wire  _T_520; // @[package.scala 32:76]
  wire  _T_522; // @[package.scala 32:76]
  wire  _T_524; // @[package.scala 32:76]
  wire [31:0] _T_525; // @[PMP.scala 62:36]
  wire [31:0] _T_527; // @[PMP.scala 62:48]
  wire [65:0] _GEN_132; // @[PMP.scala 100:53]
  wire [65:0] _T_529; // @[PMP.scala 100:53]
  wire  _T_531; // @[PMP.scala 100:78]
  wire  _T_538; // @[PMP.scala 100:78]
  wire  _T_545; // @[PMP.scala 100:78]
  wire  _T_547; // @[package.scala 32:76]
  wire  _T_549; // @[package.scala 32:76]
  wire  _T_551; // @[package.scala 32:76]
  wire  _T_552; // @[PMP.scala 100:21]
  wire  _T_565; // @[PMP.scala 109:32]
  wire [31:0] _T_585; // @[PMP.scala 113:53]
  wire [65:0] _GEN_140; // @[PMP.scala 113:40]
  wire  _T_586; // @[PMP.scala 113:40]
  wire  _T_587; // @[PMP.scala 115:21]
  wire  _T_588; // @[PMP.scala 115:62]
  wire  _T_589; // @[PMP.scala 115:41]
  wire  _T_590; // @[PMP.scala 120:58]
  wire  _T_591; // @[PMP.scala 120:8]
  wire  _T_592; // @[PMP.scala 140:10]
  wire  _T_598; // @[package.scala 32:76]
  wire  _T_600; // @[package.scala 32:76]
  wire  _T_602; // @[package.scala 32:76]
  wire [31:0] _T_603; // @[PMP.scala 62:36]
  wire [31:0] _T_605; // @[PMP.scala 62:48]
  wire [65:0] _GEN_141; // @[PMP.scala 100:53]
  wire [65:0] _T_607; // @[PMP.scala 100:53]
  wire  _T_609; // @[PMP.scala 100:78]
  wire  _T_616; // @[PMP.scala 100:78]
  wire  _T_623; // @[PMP.scala 100:78]
  wire  _T_625; // @[package.scala 32:76]
  wire  _T_627; // @[package.scala 32:76]
  wire  _T_629; // @[package.scala 32:76]
  wire  _T_630; // @[PMP.scala 100:21]
  wire  _T_643; // @[PMP.scala 109:32]
  wire [31:0] _T_663; // @[PMP.scala 113:53]
  wire [65:0] _GEN_149; // @[PMP.scala 113:40]
  wire  _T_664; // @[PMP.scala 113:40]
  wire  _T_665; // @[PMP.scala 115:21]
  wire  _T_666; // @[PMP.scala 115:62]
  wire  _T_667; // @[PMP.scala 115:41]
  wire  _T_668; // @[PMP.scala 120:58]
  wire  _T_669; // @[PMP.scala 120:8]
  wire  _T_670; // @[PMP.scala 140:10]
  wire  _T_676; // @[package.scala 32:76]
  wire  _T_678; // @[package.scala 32:76]
  wire  _T_680; // @[package.scala 32:76]
  wire [31:0] _T_681; // @[PMP.scala 62:36]
  wire [31:0] _T_683; // @[PMP.scala 62:48]
  wire [65:0] _GEN_150; // @[PMP.scala 100:53]
  wire [65:0] _T_685; // @[PMP.scala 100:53]
  wire  _T_687; // @[PMP.scala 100:78]
  wire  _T_694; // @[PMP.scala 100:78]
  wire  _T_701; // @[PMP.scala 100:78]
  wire  _T_703; // @[package.scala 32:76]
  wire  _T_705; // @[package.scala 32:76]
  wire  _T_707; // @[package.scala 32:76]
  wire  _T_708; // @[PMP.scala 100:21]
  wire  _T_721; // @[PMP.scala 109:32]
  wire [31:0] _T_741; // @[PMP.scala 113:53]
  wire [65:0] _GEN_158; // @[PMP.scala 113:40]
  wire  _T_742; // @[PMP.scala 113:40]
  wire  _T_743; // @[PMP.scala 115:21]
  wire  _T_744; // @[PMP.scala 115:62]
  wire  _T_745; // @[PMP.scala 115:41]
  wire  _T_746; // @[PMP.scala 120:58]
  wire  _T_747; // @[PMP.scala 120:8]
  wire  _T_748; // @[PMP.scala 140:10]
  wire  _T_754; // @[package.scala 32:76]
  wire  _T_756; // @[package.scala 32:76]
  wire  _T_758; // @[package.scala 32:76]
  wire [31:0] _T_759; // @[PMP.scala 62:36]
  wire [31:0] _T_761; // @[PMP.scala 62:48]
  wire [65:0] _GEN_159; // @[PMP.scala 100:53]
  wire [65:0] _T_763; // @[PMP.scala 100:53]
  wire  _T_765; // @[PMP.scala 100:78]
  wire  _T_772; // @[PMP.scala 100:78]
  wire  _T_779; // @[PMP.scala 100:78]
  wire  _T_781; // @[package.scala 32:76]
  wire  _T_783; // @[package.scala 32:76]
  wire  _T_785; // @[package.scala 32:76]
  wire  _T_786; // @[PMP.scala 100:21]
  wire  _T_799; // @[PMP.scala 109:32]
  wire [31:0] _T_819; // @[PMP.scala 113:53]
  wire [65:0] _GEN_167; // @[PMP.scala 113:40]
  wire  _T_820; // @[PMP.scala 113:40]
  wire  _T_821; // @[PMP.scala 115:21]
  wire  _T_822; // @[PMP.scala 115:62]
  wire  _T_823; // @[PMP.scala 115:41]
  wire  _T_824; // @[PMP.scala 120:58]
  wire  _T_825; // @[PMP.scala 120:8]
  wire  _T_826; // @[PMP.scala 140:10]
  wire  _T_832; // @[package.scala 32:76]
  wire  _T_834; // @[package.scala 32:76]
  wire  _T_836; // @[package.scala 32:76]
  wire [31:0] _T_837; // @[PMP.scala 62:36]
  wire [31:0] _T_839; // @[PMP.scala 62:48]
  wire [65:0] _GEN_168; // @[PMP.scala 100:53]
  wire [65:0] _T_841; // @[PMP.scala 100:53]
  wire  _T_843; // @[PMP.scala 100:78]
  wire  _T_850; // @[PMP.scala 100:78]
  wire  _T_857; // @[PMP.scala 100:78]
  wire  _T_859; // @[package.scala 32:76]
  wire  _T_861; // @[package.scala 32:76]
  wire  _T_863; // @[package.scala 32:76]
  wire  _T_864; // @[PMP.scala 100:21]
  wire  _T_877; // @[PMP.scala 109:32]
  wire [31:0] _T_897; // @[PMP.scala 113:53]
  wire [65:0] _GEN_176; // @[PMP.scala 113:40]
  wire  _T_898; // @[PMP.scala 113:40]
  wire  _T_899; // @[PMP.scala 115:21]
  wire  _T_900; // @[PMP.scala 115:62]
  wire  _T_901; // @[PMP.scala 115:41]
  wire  _T_902; // @[PMP.scala 120:58]
  wire  _T_903; // @[PMP.scala 120:8]
  wire  _T_904; // @[PMP.scala 140:10]
  wire  _T_910; // @[package.scala 32:76]
  wire  _T_912; // @[package.scala 32:76]
  wire  _T_914; // @[package.scala 32:76]
  wire [31:0] _T_915; // @[PMP.scala 62:36]
  wire [31:0] _T_917; // @[PMP.scala 62:48]
  wire [65:0] _GEN_177; // @[PMP.scala 100:53]
  wire [65:0] _T_919; // @[PMP.scala 100:53]
  wire  _T_921; // @[PMP.scala 100:78]
  wire  _T_928; // @[PMP.scala 100:78]
  wire  _T_935; // @[PMP.scala 100:78]
  wire  _T_937; // @[package.scala 32:76]
  wire  _T_939; // @[package.scala 32:76]
  wire  _T_941; // @[package.scala 32:76]
  wire  _T_942; // @[PMP.scala 100:21]
  wire  _T_955; // @[PMP.scala 109:32]
  wire [31:0] _T_975; // @[PMP.scala 113:53]
  wire [65:0] _GEN_185; // @[PMP.scala 113:40]
  wire  _T_976; // @[PMP.scala 113:40]
  wire  _T_977; // @[PMP.scala 115:21]
  wire  _T_978; // @[PMP.scala 115:62]
  wire  _T_979; // @[PMP.scala 115:41]
  wire  _T_980; // @[PMP.scala 120:58]
  wire  _T_981; // @[PMP.scala 120:8]
  wire  pmpHomogeneous; // @[PMP.scala 140:10]
  wire  homogeneous; // @[PTW.scala 269:36]
  wire  _T_986; // @[Conditional.scala 37:30]
  wire [2:0] _T_988; // @[PTW.scala 291:26]
  wire [2:0] _GEN_40; // @[PTW.scala 290:32]
  wire  _T_990; // @[PTW.scala 293:39]
  wire  _T_991; // @[Conditional.scala 37:30]
  wire [1:0] _T_993; // @[PTW.scala 297:24]
  wire [2:0] _T_994; // @[PTW.scala 299:26]
  wire [2:0] _GEN_42; // @[PTW.scala 296:28]
  wire  _T_995; // @[Conditional.scala 37:30]
  wire  _T_997; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_46; // @[PTW.scala 308:35]
  wire  _GEN_47; // @[PTW.scala 308:35]
  wire  _GEN_48; // @[PTW.scala 308:35]
  wire  _T_1000; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_54; // @[Conditional.scala 39:67]
  wire  _GEN_55; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_59; // @[Conditional.scala 39:67]
  wire  _GEN_60; // @[Conditional.scala 39:67]
  wire  _GEN_61; // @[Conditional.scala 39:67]
  wire  _GEN_62; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_65; // @[Conditional.scala 39:67]
  wire  _GEN_67; // @[Conditional.scala 39:67]
  wire  _GEN_68; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_72; // @[Conditional.scala 39:67]
  wire  _GEN_74; // @[Conditional.scala 39:67]
  wire  _GEN_75; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_77; // @[Conditional.scala 40:58]
  wire  _GEN_80; // @[Conditional.scala 40:58]
  wire  _GEN_81; // @[Conditional.scala 40:58]
  wire  _T_1006; // @[PTW.scala 333:15]
  wire  _T_1008; // @[PTW.scala 333:40]
  wire  _T_1010; // @[PTW.scala 334:25]
  wire [53:0] pte_2_ppn; // @[PTW.scala 327:13]
  wire [53:0] _T_1012_ppn; // @[PTW.scala 335:8]
  wire [53:0] pte_1_ppn; // @[PTW.scala 327:13]
  wire [53:0] _T_1013_ppn; // @[PTW.scala 334:8]
  wire  _T_1013_d; // @[PTW.scala 334:8]
  wire  _T_1013_a; // @[PTW.scala 334:8]
  wire  _T_1013_g; // @[PTW.scala 334:8]
  wire  _T_1013_u; // @[PTW.scala 334:8]
  wire  _T_1013_x; // @[PTW.scala 334:8]
  wire  _T_1013_w; // @[PTW.scala 334:8]
  wire  _T_1013_r; // @[PTW.scala 334:8]
  wire  _T_1013_v; // @[PTW.scala 334:8]
  wire [53:0] _T_1014_ppn; // @[PTW.scala 333:8]
  wire  _T_1014_d; // @[PTW.scala 333:8]
  wire  _T_1014_a; // @[PTW.scala 333:8]
  wire  _T_1014_g; // @[PTW.scala 333:8]
  wire  _T_1014_u; // @[PTW.scala 333:8]
  wire  _T_1014_x; // @[PTW.scala 333:8]
  wire  _T_1014_w; // @[PTW.scala 333:8]
  wire  _T_1014_r; // @[PTW.scala 333:8]
  wire  _T_1014_v; // @[PTW.scala 333:8]
  wire  _GEN_83; // @[PTW.scala 341:28]
  wire  _GEN_84; // @[PTW.scala 341:28]
  wire  _T_1027; // @[PTW.scala 346:18]
  wire  _T_1029; // @[PTW.scala 346:11]
  wire  ae; // @[PTW.scala 352:22]
  wire [2:0] _GEN_95; // @[PTW.scala 347:21]
  wire [2:0] _GEN_101; // @[PTW.scala 345:25]
  wire  _T_1043; // @[PTW.scala 363:18]
  wire  _T_1045; // @[PTW.scala 363:11]
  reg [19:0] PTW_state; // @[Register tracking PTW state]
  reg [31:0] _RAND_37;
  reg  PTW_cov [0:1048575]; // @[Coverage map for PTW]
  reg [31:0] _RAND_38;
  wire  PTW_cov_read_data; // @[Coverage map for PTW]
  wire [19:0] PTW_cov_read_addr; // @[Coverage map for PTW]
  wire  PTW_cov_write_data; // @[Coverage map for PTW]
  wire [19:0] PTW_cov_write_addr; // @[Coverage map for PTW]
  wire  PTW_cov_write_mask; // @[Coverage map for PTW]
  wire  PTW_cov_write_en; // @[Coverage map for PTW]
  reg [29:0] PTW_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_39;
  wire [10:0] valid_shl;
  wire [19:0] valid_pad;
  wire [11:0] invalidated_shl;
  wire [19:0] invalidated_pad;
  wire [12:0] state_shl;
  wire [19:0] state_pad;
  wire [6:0] _T_56_shl;
  wire [19:0] _T_56_pad;
  wire [15:0] count_shl;
  wire [19:0] count_pad;
  wire [1:0] mem_resp_valid_shl;
  wire [19:0] mem_resp_valid_pad;
  wire [19:0] PTW_xor4;
  wire [19:0] PTW_xor1;
  wire [19:0] PTW_xor6;
  wire [19:0] PTW_xor2;
  wire [19:0] PTW_xor0;
  wire [29:0] arb_sum;
  wire [29:0] OptimizationBarrier_sum;
  wire [29:0] OptimizationBarrier_1_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  arb_metaAssert_wire;
  wire  OptimizationBarrier_metaAssert_wire;
  wire  OptimizationBarrier_1_metaAssert_wire;
  wire  PTW_or1;
  wire  PTW_or6;
  wire  PTW_or2;
  wire  PTW_or0;
  reg  PTW_metaAssert;
  reg [31:0] _RAND_40;
  Arbiter arb ( // @[PTW.scala 105:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_bits_addr(arb_io_in_0_bits_bits_addr),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_valid(arb_io_in_1_bits_valid),
    .io_in_1_bits_bits_addr(arb_io_in_1_bits_bits_addr),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_valid(arb_io_out_bits_valid),
    .io_out_bits_bits_addr(arb_io_out_bits_bits_addr),
    .io_chosen(arb_io_chosen),
    .io_covSum(arb_io_covSum),
    .metaAssert(arb_metaAssert)
  );
  OptimizationBarrier_117 OptimizationBarrier ( // @[package.scala 236:25]
    .io_x(OptimizationBarrier_io_x),
    .io_y(OptimizationBarrier_io_y),
    .io_covSum(OptimizationBarrier_io_covSum),
    .metaAssert(OptimizationBarrier_metaAssert)
  );
  OptimizationBarrier_118 OptimizationBarrier_1 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_1_io_x_ppn),
    .io_x_d(OptimizationBarrier_1_io_x_d),
    .io_x_a(OptimizationBarrier_1_io_x_a),
    .io_x_g(OptimizationBarrier_1_io_x_g),
    .io_x_u(OptimizationBarrier_1_io_x_u),
    .io_x_x(OptimizationBarrier_1_io_x_x),
    .io_x_w(OptimizationBarrier_1_io_x_w),
    .io_x_r(OptimizationBarrier_1_io_x_r),
    .io_x_v(OptimizationBarrier_1_io_x_v),
    .io_y_ppn(OptimizationBarrier_1_io_y_ppn),
    .io_y_d(OptimizationBarrier_1_io_y_d),
    .io_y_a(OptimizationBarrier_1_io_y_a),
    .io_y_g(OptimizationBarrier_1_io_y_g),
    .io_y_u(OptimizationBarrier_1_io_y_u),
    .io_y_x(OptimizationBarrier_1_io_y_x),
    .io_y_w(OptimizationBarrier_1_io_y_w),
    .io_y_r(OptimizationBarrier_1_io_y_r),
    .io_y_v(OptimizationBarrier_1_io_y_v),
    .io_covSum(OptimizationBarrier_1_io_covSum),
    .metaAssert(OptimizationBarrier_1_metaAssert)
  );
  assign _T_2 = state != 3'h0; // @[PTW.scala 111:24]
  assign tmp_v = mem_resp_data[0]; // @[PTW.scala 139:33]
  assign tmp_r = mem_resp_data[1]; // @[PTW.scala 139:33]
  assign tmp_w = mem_resp_data[2]; // @[PTW.scala 139:33]
  assign tmp_x = mem_resp_data[3]; // @[PTW.scala 139:33]
  assign tmp_u = mem_resp_data[4]; // @[PTW.scala 139:33]
  assign tmp_g = mem_resp_data[5]; // @[PTW.scala 139:33]
  assign tmp_a = mem_resp_data[6]; // @[PTW.scala 139:33]
  assign tmp_d = mem_resp_data[7]; // @[PTW.scala 139:33]
  assign tmp_ppn = mem_resp_data[63:10]; // @[PTW.scala 139:33]
  assign _T_19 = tmp_r | tmp_w; // @[PTW.scala 142:17]
  assign _T_20 = _T_19 | tmp_x; // @[PTW.scala 142:26]
  assign _T_21 = count <= 2'h0; // @[PTW.scala 145:21]
  assign _T_23 = tmp_ppn[17:9] != 9'h0; // @[PTW.scala 145:95]
  assign _T_24 = _T_21 & _T_23; // @[PTW.scala 145:26]
  assign _GEN_0 = _T_24 ? 1'h0 : tmp_v; // @[PTW.scala 145:102]
  assign _T_25 = count <= 2'h1; // @[PTW.scala 145:21]
  assign _T_27 = tmp_ppn[8:0] != 9'h0; // @[PTW.scala 145:95]
  assign _T_28 = _T_25 & _T_27; // @[PTW.scala 145:26]
  assign _GEN_1 = _T_28 ? 1'h0 : _GEN_0; // @[PTW.scala 145:102]
  assign res_v = _T_20 ? _GEN_1 : tmp_v; // @[PTW.scala 142:36]
  assign invalid_paddr = tmp_ppn[53:20] != 34'h0; // @[PTW.scala 147:32]
  assign _T_31 = res_v & ~tmp_r; // @[PTW.scala 68:33]
  assign _T_33 = _T_31 & ~tmp_w; // @[PTW.scala 68:39]
  assign _T_35 = _T_33 & ~tmp_x; // @[PTW.scala 68:45]
  assign _T_37 = _T_35 & ~invalid_paddr; // @[PTW.scala 149:30]
  assign _T_38 = count < 2'h2; // @[PTW.scala 149:57]
  assign traverse = _T_37 & _T_38; // @[PTW.scala 149:48]
  assign vpn_idxs_0 = r_req_addr[26:18]; // @[PTW.scala 151:60]
  assign vpn_idxs_1 = r_req_addr[17:9]; // @[PTW.scala 151:90]
  assign vpn_idxs_2 = r_req_addr[8:0]; // @[PTW.scala 151:90]
  assign _T_42 = count == 2'h1; // @[package.scala 32:86]
  assign _T_43 = _T_42 ? vpn_idxs_1 : vpn_idxs_0; // @[package.scala 32:76]
  assign _T_44 = count == 2'h2; // @[package.scala 32:86]
  assign _T_45 = _T_44 ? vpn_idxs_2 : _T_43; // @[package.scala 32:76]
  assign _T_46 = count == 2'h3; // @[package.scala 32:86]
  assign vpn_idx = _T_46 ? vpn_idxs_2 : _T_45; // @[package.scala 32:76]
  assign _T_47 = {r_pte_ppn,vpn_idx}; // @[Cat.scala 29:58]
  assign pte_addr = {_T_47, 3'h0}; // @[PTW.scala 153:29]
  assign choices_0 = {r_pte_ppn[53:18],r_req_addr[17:0]}; // @[Cat.scala 29:58]
  assign choices_1 = {r_pte_ppn[53:9],vpn_idxs_2}; // @[Cat.scala 29:58]
  assign fragmented_superpage_ppn = count[0] ? choices_1 : choices_0; // @[package.scala 32:76]
  assign _T_55 = arb_io_out_ready & arb_io_out_valid; // @[Decoupled.scala 40:37]
  assign _GEN_108 = {{34'd0}, tags_0}; // @[PTW.scala 172:27]
  assign _T_57 = _GEN_108 == pte_addr; // @[PTW.scala 172:27]
  assign _GEN_109 = {{34'd0}, tags_1}; // @[PTW.scala 172:27]
  assign _T_58 = _GEN_109 == pte_addr; // @[PTW.scala 172:27]
  assign _GEN_110 = {{34'd0}, tags_2}; // @[PTW.scala 172:27]
  assign _T_59 = _GEN_110 == pte_addr; // @[PTW.scala 172:27]
  assign _GEN_111 = {{34'd0}, tags_3}; // @[PTW.scala 172:27]
  assign _T_60 = _GEN_111 == pte_addr; // @[PTW.scala 172:27]
  assign _GEN_112 = {{34'd0}, tags_4}; // @[PTW.scala 172:27]
  assign _T_61 = _GEN_112 == pte_addr; // @[PTW.scala 172:27]
  assign _GEN_113 = {{34'd0}, tags_5}; // @[PTW.scala 172:27]
  assign _T_62 = _GEN_113 == pte_addr; // @[PTW.scala 172:27]
  assign _GEN_114 = {{34'd0}, tags_6}; // @[PTW.scala 172:27]
  assign _T_63 = _GEN_114 == pte_addr; // @[PTW.scala 172:27]
  assign _GEN_115 = {{34'd0}, tags_7}; // @[PTW.scala 172:27]
  assign _T_64 = _GEN_115 == pte_addr; // @[PTW.scala 172:27]
  assign _T_71 = {_T_64,_T_63,_T_62,_T_61,_T_60,_T_59,_T_58,_T_57}; // @[Cat.scala 29:58]
  assign hits = _T_71 & valid; // @[PTW.scala 172:48]
  assign hit = |hits; // @[PTW.scala 173:20]
  assign _T_72 = mem_resp_valid & traverse; // @[PTW.scala 174:26]
  assign _T_74 = _T_72 & ~hit; // @[PTW.scala 174:38]
  assign _T_76 = _T_74 & ~invalidated; // @[PTW.scala 174:46]
  assign _T_77 = &valid; // @[PTW.scala 175:25]
  assign _T_86 = _T_56[5] ? _T_56[4] : _T_56[3]; // @[Replacement.scala 240:16]
  assign _T_87 = {_T_56[5],_T_86}; // @[Cat.scala 29:58]
  assign _T_93 = _T_56[2] ? _T_56[1] : _T_56[0]; // @[Replacement.scala 240:16]
  assign _T_94 = {_T_56[2],_T_93}; // @[Cat.scala 29:58]
  assign _T_95 = _T_56[6] ? _T_87 : _T_94; // @[Replacement.scala 240:16]
  assign _T_96 = {_T_56[6],_T_95}; // @[Cat.scala 29:58]
  assign _T_98 = ~valid[0]; // @[OneHot.scala 47:40]
  assign _T_99 = ~valid[1]; // @[OneHot.scala 47:40]
  assign _T_100 = ~valid[2]; // @[OneHot.scala 47:40]
  assign _T_101 = ~valid[3]; // @[OneHot.scala 47:40]
  assign _T_102 = ~valid[4]; // @[OneHot.scala 47:40]
  assign _T_103 = ~valid[5]; // @[OneHot.scala 47:40]
  assign _T_104 = ~valid[6]; // @[OneHot.scala 47:40]
  assign _T_106 = _T_104 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  assign _T_107 = _T_103 ? 3'h5 : _T_106; // @[Mux.scala 47:69]
  assign _T_108 = _T_102 ? 3'h4 : _T_107; // @[Mux.scala 47:69]
  assign _T_109 = _T_101 ? 3'h3 : _T_108; // @[Mux.scala 47:69]
  assign _T_110 = _T_100 ? 3'h2 : _T_109; // @[Mux.scala 47:69]
  assign _T_111 = _T_99 ? 3'h1 : _T_110; // @[Mux.scala 47:69]
  assign _T_112 = _T_98 ? 3'h0 : _T_111; // @[Mux.scala 47:69]
  assign r = _T_77 ? _T_96 : _T_112; // @[PTW.scala 175:18]
  assign _T_113 = 8'h1 << r; // @[OneHot.scala 58:35]
  assign _T_114 = valid | _T_113; // @[PTW.scala 176:22]
  assign res_ppn = {{34'd0}, tmp_ppn[19:0]}; // @[PTW.scala 141:13]
  assign _T_115 = state == 3'h1; // @[PTW.scala 180:24]
  assign _T_116 = hit & _T_115; // @[PTW.scala 180:15]
  assign _T_119 = |hits[7:4]; // @[OneHot.scala 32:14]
  assign _T_120 = hits[7:4] | hits[3:0]; // @[OneHot.scala 32:28]
  assign _T_123 = |_T_120[3:2]; // @[OneHot.scala 32:14]
  assign _T_124 = _T_120[3:2] | _T_120[1:0]; // @[OneHot.scala 32:28]
  assign _T_127 = {_T_119,_T_123,_T_124[1]}; // @[Cat.scala 29:58]
  assign _T_141 = _T_127[1] ? ~_T_127[0] : _T_56[4]; // @[Replacement.scala 193:16]
  assign _T_145 = _T_127[1] ? _T_56[3] : ~_T_127[0]; // @[Replacement.scala 196:16]
  assign _T_147 = {~_T_127[1],_T_141,_T_145}; // @[Cat.scala 29:58]
  assign _T_148 = _T_127[2] ? _T_147 : _T_56[5:3]; // @[Replacement.scala 193:16]
  assign _T_157 = _T_127[1] ? ~_T_127[0] : _T_56[1]; // @[Replacement.scala 193:16]
  assign _T_161 = _T_127[1] ? _T_56[0] : ~_T_127[0]; // @[Replacement.scala 196:16]
  assign _T_163 = {~_T_127[1],_T_157,_T_161}; // @[Cat.scala 29:58]
  assign _T_164 = _T_127[2] ? _T_56[2:0] : _T_163; // @[Replacement.scala 196:16]
  assign _T_166 = {~_T_127[2],_T_148,_T_164}; // @[Cat.scala 29:58]
  assign _T_168 = io_dpath_sfence_valid & ~io_dpath_sfence_bits_rs1; // @[PTW.scala 181:33]
  assign pte_cache_hit = hit & _T_38; // @[PTW.scala 186:10]
  assign _T_186 = hits[0] ? data_0 : 20'h0; // @[Mux.scala 27:72]
  assign _T_187 = hits[1] ? data_1 : 20'h0; // @[Mux.scala 27:72]
  assign _T_188 = hits[2] ? data_2 : 20'h0; // @[Mux.scala 27:72]
  assign _T_189 = hits[3] ? data_3 : 20'h0; // @[Mux.scala 27:72]
  assign _T_190 = hits[4] ? data_4 : 20'h0; // @[Mux.scala 27:72]
  assign _T_191 = hits[5] ? data_5 : 20'h0; // @[Mux.scala 27:72]
  assign _T_192 = hits[6] ? data_6 : 20'h0; // @[Mux.scala 27:72]
  assign _T_193 = hits[7] ? data_7 : 20'h0; // @[Mux.scala 27:72]
  assign _T_194 = _T_186 | _T_187; // @[Mux.scala 27:72]
  assign _T_195 = _T_194 | _T_188; // @[Mux.scala 27:72]
  assign _T_196 = _T_195 | _T_189; // @[Mux.scala 27:72]
  assign _T_197 = _T_196 | _T_190; // @[Mux.scala 27:72]
  assign _T_198 = _T_197 | _T_191; // @[Mux.scala 27:72]
  assign _T_199 = _T_198 | _T_192; // @[Mux.scala 27:72]
  assign pte_cache_data = _T_199 | _T_193; // @[Mux.scala 27:72]
  assign _T_202 = invalidated & _T_2; // @[PTW.scala 245:56]
  assign _T_205 = state == 3'h3; // @[PTW.scala 247:48]
  assign _T_215 = pte_addr ^ 66'hc000000; // @[Parameters.scala 137:31]
  assign _T_216 = {1'b0,$signed(_T_215)}; // @[Parameters.scala 137:49]
  assign _T_218 = $signed(_T_216) & -67'sh4000000; // @[Parameters.scala 137:52]
  assign _T_219 = $signed(_T_218) == 67'sh0; // @[Parameters.scala 137:67]
  assign _T_220 = pte_addr ^ 66'h60000000; // @[Parameters.scala 137:31]
  assign _T_221 = {1'b0,$signed(_T_220)}; // @[Parameters.scala 137:49]
  assign _T_223 = $signed(_T_221) & -67'sh20000000; // @[Parameters.scala 137:52]
  assign _T_224 = $signed(_T_223) == 67'sh0; // @[Parameters.scala 137:67]
  assign _T_225 = pte_addr ^ 66'h80000000; // @[Parameters.scala 137:31]
  assign _T_226 = {1'b0,$signed(_T_225)}; // @[Parameters.scala 137:49]
  assign _T_228 = $signed(_T_226) & -67'sh10000000; // @[Parameters.scala 137:52]
  assign _T_229 = $signed(_T_228) == 67'sh0; // @[Parameters.scala 137:67]
  assign _T_231 = _T_219 | _T_224; // @[TLBPermissions.scala 98:65]
  assign pmaPgLevelHomogeneous_1 = _T_231 | _T_229; // @[TLBPermissions.scala 98:65]
  assign _T_235 = {1'b0,$signed(pte_addr)}; // @[Parameters.scala 137:49]
  assign _T_262 = $signed(_T_235) & -67'sh1000; // @[Parameters.scala 137:52]
  assign _T_263 = $signed(_T_262) == 67'sh0; // @[Parameters.scala 137:67]
  assign _T_264 = pte_addr ^ 66'h3000; // @[Parameters.scala 137:31]
  assign _T_265 = {1'b0,$signed(_T_264)}; // @[Parameters.scala 137:49]
  assign _T_267 = $signed(_T_265) & -67'sh1000; // @[Parameters.scala 137:52]
  assign _T_268 = $signed(_T_267) == 67'sh0; // @[Parameters.scala 137:67]
  assign _T_269 = pte_addr ^ 66'h10000; // @[Parameters.scala 137:31]
  assign _T_270 = {1'b0,$signed(_T_269)}; // @[Parameters.scala 137:49]
  assign _T_272 = $signed(_T_270) & -67'sh10000; // @[Parameters.scala 137:52]
  assign _T_273 = $signed(_T_272) == 67'sh0; // @[Parameters.scala 137:67]
  assign _T_274 = pte_addr ^ 66'h2000000; // @[Parameters.scala 137:31]
  assign _T_275 = {1'b0,$signed(_T_274)}; // @[Parameters.scala 137:49]
  assign _T_277 = $signed(_T_275) & -67'sh10000; // @[Parameters.scala 137:52]
  assign _T_278 = $signed(_T_277) == 67'sh0; // @[Parameters.scala 137:67]
  assign _T_295 = _T_263 | _T_268; // @[TLBPermissions.scala 98:65]
  assign _T_296 = _T_295 | _T_273; // @[TLBPermissions.scala 98:65]
  assign _T_297 = _T_296 | _T_278; // @[TLBPermissions.scala 98:65]
  assign _T_298 = _T_297 | _T_219; // @[TLBPermissions.scala 98:65]
  assign _T_299 = _T_298 | _T_224; // @[TLBPermissions.scala 98:65]
  assign pmaPgLevelHomogeneous_2 = _T_299 | _T_229; // @[TLBPermissions.scala 98:65]
  assign _T_352 = _T_42 & pmaPgLevelHomogeneous_1; // @[package.scala 32:76]
  assign _T_354 = _T_44 ? pmaPgLevelHomogeneous_2 : _T_352; // @[package.scala 32:76]
  assign pmaHomogeneous = _T_46 ? pmaPgLevelHomogeneous_2 : _T_354; // @[package.scala 32:76]
  assign _T_357 = {pte_addr[65:12], 12'h0}; // @[PTW.scala 268:92]
  assign _T_364 = _T_42 ? io_dpath_pmp_0_mask[20] : io_dpath_pmp_0_mask[29]; // @[package.scala 32:76]
  assign _T_366 = _T_44 ? io_dpath_pmp_0_mask[11] : _T_364; // @[package.scala 32:76]
  assign _T_368 = _T_46 ? io_dpath_pmp_0_mask[11] : _T_366; // @[package.scala 32:76]
  assign _T_369 = {io_dpath_pmp_0_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_371 = ~_T_369 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_116 = {{34'd0}, ~_T_371}; // @[PMP.scala 100:53]
  assign _T_373 = _T_357 ^ _GEN_116; // @[PMP.scala 100:53]
  assign _T_375 = _T_373[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _T_382 = _T_373[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _T_389 = _T_373[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _T_391 = _T_42 ? _T_382 : _T_375; // @[package.scala 32:76]
  assign _T_393 = _T_44 ? _T_389 : _T_391; // @[package.scala 32:76]
  assign _T_395 = _T_46 ? _T_389 : _T_393; // @[package.scala 32:76]
  assign _T_396 = _T_368 | _T_395; // @[PMP.scala 100:21]
  assign _T_409 = _T_357 < _GEN_116; // @[PMP.scala 109:32]
  assign _T_412 = _T_42 ? 32'hffe00000 : 32'hc0000000; // @[package.scala 32:76]
  assign _T_414 = _T_44 ? 32'hfffff000 : _T_412; // @[package.scala 32:76]
  assign _T_416 = _T_46 ? 32'hfffff000 : _T_414; // @[package.scala 32:76]
  assign _GEN_120 = {{34'd0}, _T_416}; // @[PMP.scala 112:30]
  assign _T_417 = _T_357 & _GEN_120; // @[PMP.scala 112:30]
  assign _T_429 = ~_T_371 & _T_416; // @[PMP.scala 113:53]
  assign _GEN_122 = {{34'd0}, _T_429}; // @[PMP.scala 113:40]
  assign _T_430 = _T_417 < _GEN_122; // @[PMP.scala 113:40]
  assign _T_433 = ~_T_409 | _T_430; // @[PMP.scala 115:41]
  assign _T_434 = ~io_dpath_pmp_0_cfg_a[0] | _T_433; // @[PMP.scala 120:58]
  assign _T_435 = io_dpath_pmp_0_cfg_a[1] ? _T_396 : _T_434; // @[PMP.scala 120:8]
  assign _T_442 = _T_42 ? io_dpath_pmp_1_mask[20] : io_dpath_pmp_1_mask[29]; // @[package.scala 32:76]
  assign _T_444 = _T_44 ? io_dpath_pmp_1_mask[11] : _T_442; // @[package.scala 32:76]
  assign _T_446 = _T_46 ? io_dpath_pmp_1_mask[11] : _T_444; // @[package.scala 32:76]
  assign _T_447 = {io_dpath_pmp_1_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_449 = ~_T_447 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_123 = {{34'd0}, ~_T_449}; // @[PMP.scala 100:53]
  assign _T_451 = _T_357 ^ _GEN_123; // @[PMP.scala 100:53]
  assign _T_453 = _T_451[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _T_460 = _T_451[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _T_467 = _T_451[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _T_469 = _T_42 ? _T_460 : _T_453; // @[package.scala 32:76]
  assign _T_471 = _T_44 ? _T_467 : _T_469; // @[package.scala 32:76]
  assign _T_473 = _T_46 ? _T_467 : _T_471; // @[package.scala 32:76]
  assign _T_474 = _T_446 | _T_473; // @[PMP.scala 100:21]
  assign _T_487 = _T_357 < _GEN_123; // @[PMP.scala 109:32]
  assign _T_507 = ~_T_449 & _T_416; // @[PMP.scala 113:53]
  assign _GEN_131 = {{34'd0}, _T_507}; // @[PMP.scala 113:40]
  assign _T_508 = _T_417 < _GEN_131; // @[PMP.scala 113:40]
  assign _T_509 = _T_430 | ~_T_487; // @[PMP.scala 115:21]
  assign _T_510 = ~_T_409 & _T_508; // @[PMP.scala 115:62]
  assign _T_511 = _T_509 | _T_510; // @[PMP.scala 115:41]
  assign _T_512 = ~io_dpath_pmp_1_cfg_a[0] | _T_511; // @[PMP.scala 120:58]
  assign _T_513 = io_dpath_pmp_1_cfg_a[1] ? _T_474 : _T_512; // @[PMP.scala 120:8]
  assign _T_514 = _T_435 & _T_513; // @[PMP.scala 140:10]
  assign _T_520 = _T_42 ? io_dpath_pmp_2_mask[20] : io_dpath_pmp_2_mask[29]; // @[package.scala 32:76]
  assign _T_522 = _T_44 ? io_dpath_pmp_2_mask[11] : _T_520; // @[package.scala 32:76]
  assign _T_524 = _T_46 ? io_dpath_pmp_2_mask[11] : _T_522; // @[package.scala 32:76]
  assign _T_525 = {io_dpath_pmp_2_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_527 = ~_T_525 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_132 = {{34'd0}, ~_T_527}; // @[PMP.scala 100:53]
  assign _T_529 = _T_357 ^ _GEN_132; // @[PMP.scala 100:53]
  assign _T_531 = _T_529[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _T_538 = _T_529[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _T_545 = _T_529[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _T_547 = _T_42 ? _T_538 : _T_531; // @[package.scala 32:76]
  assign _T_549 = _T_44 ? _T_545 : _T_547; // @[package.scala 32:76]
  assign _T_551 = _T_46 ? _T_545 : _T_549; // @[package.scala 32:76]
  assign _T_552 = _T_524 | _T_551; // @[PMP.scala 100:21]
  assign _T_565 = _T_357 < _GEN_132; // @[PMP.scala 109:32]
  assign _T_585 = ~_T_527 & _T_416; // @[PMP.scala 113:53]
  assign _GEN_140 = {{34'd0}, _T_585}; // @[PMP.scala 113:40]
  assign _T_586 = _T_417 < _GEN_140; // @[PMP.scala 113:40]
  assign _T_587 = _T_508 | ~_T_565; // @[PMP.scala 115:21]
  assign _T_588 = ~_T_487 & _T_586; // @[PMP.scala 115:62]
  assign _T_589 = _T_587 | _T_588; // @[PMP.scala 115:41]
  assign _T_590 = ~io_dpath_pmp_2_cfg_a[0] | _T_589; // @[PMP.scala 120:58]
  assign _T_591 = io_dpath_pmp_2_cfg_a[1] ? _T_552 : _T_590; // @[PMP.scala 120:8]
  assign _T_592 = _T_514 & _T_591; // @[PMP.scala 140:10]
  assign _T_598 = _T_42 ? io_dpath_pmp_3_mask[20] : io_dpath_pmp_3_mask[29]; // @[package.scala 32:76]
  assign _T_600 = _T_44 ? io_dpath_pmp_3_mask[11] : _T_598; // @[package.scala 32:76]
  assign _T_602 = _T_46 ? io_dpath_pmp_3_mask[11] : _T_600; // @[package.scala 32:76]
  assign _T_603 = {io_dpath_pmp_3_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_605 = ~_T_603 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_141 = {{34'd0}, ~_T_605}; // @[PMP.scala 100:53]
  assign _T_607 = _T_357 ^ _GEN_141; // @[PMP.scala 100:53]
  assign _T_609 = _T_607[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _T_616 = _T_607[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _T_623 = _T_607[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _T_625 = _T_42 ? _T_616 : _T_609; // @[package.scala 32:76]
  assign _T_627 = _T_44 ? _T_623 : _T_625; // @[package.scala 32:76]
  assign _T_629 = _T_46 ? _T_623 : _T_627; // @[package.scala 32:76]
  assign _T_630 = _T_602 | _T_629; // @[PMP.scala 100:21]
  assign _T_643 = _T_357 < _GEN_141; // @[PMP.scala 109:32]
  assign _T_663 = ~_T_605 & _T_416; // @[PMP.scala 113:53]
  assign _GEN_149 = {{34'd0}, _T_663}; // @[PMP.scala 113:40]
  assign _T_664 = _T_417 < _GEN_149; // @[PMP.scala 113:40]
  assign _T_665 = _T_586 | ~_T_643; // @[PMP.scala 115:21]
  assign _T_666 = ~_T_565 & _T_664; // @[PMP.scala 115:62]
  assign _T_667 = _T_665 | _T_666; // @[PMP.scala 115:41]
  assign _T_668 = ~io_dpath_pmp_3_cfg_a[0] | _T_667; // @[PMP.scala 120:58]
  assign _T_669 = io_dpath_pmp_3_cfg_a[1] ? _T_630 : _T_668; // @[PMP.scala 120:8]
  assign _T_670 = _T_592 & _T_669; // @[PMP.scala 140:10]
  assign _T_676 = _T_42 ? io_dpath_pmp_4_mask[20] : io_dpath_pmp_4_mask[29]; // @[package.scala 32:76]
  assign _T_678 = _T_44 ? io_dpath_pmp_4_mask[11] : _T_676; // @[package.scala 32:76]
  assign _T_680 = _T_46 ? io_dpath_pmp_4_mask[11] : _T_678; // @[package.scala 32:76]
  assign _T_681 = {io_dpath_pmp_4_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_683 = ~_T_681 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_150 = {{34'd0}, ~_T_683}; // @[PMP.scala 100:53]
  assign _T_685 = _T_357 ^ _GEN_150; // @[PMP.scala 100:53]
  assign _T_687 = _T_685[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _T_694 = _T_685[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _T_701 = _T_685[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _T_703 = _T_42 ? _T_694 : _T_687; // @[package.scala 32:76]
  assign _T_705 = _T_44 ? _T_701 : _T_703; // @[package.scala 32:76]
  assign _T_707 = _T_46 ? _T_701 : _T_705; // @[package.scala 32:76]
  assign _T_708 = _T_680 | _T_707; // @[PMP.scala 100:21]
  assign _T_721 = _T_357 < _GEN_150; // @[PMP.scala 109:32]
  assign _T_741 = ~_T_683 & _T_416; // @[PMP.scala 113:53]
  assign _GEN_158 = {{34'd0}, _T_741}; // @[PMP.scala 113:40]
  assign _T_742 = _T_417 < _GEN_158; // @[PMP.scala 113:40]
  assign _T_743 = _T_664 | ~_T_721; // @[PMP.scala 115:21]
  assign _T_744 = ~_T_643 & _T_742; // @[PMP.scala 115:62]
  assign _T_745 = _T_743 | _T_744; // @[PMP.scala 115:41]
  assign _T_746 = ~io_dpath_pmp_4_cfg_a[0] | _T_745; // @[PMP.scala 120:58]
  assign _T_747 = io_dpath_pmp_4_cfg_a[1] ? _T_708 : _T_746; // @[PMP.scala 120:8]
  assign _T_748 = _T_670 & _T_747; // @[PMP.scala 140:10]
  assign _T_754 = _T_42 ? io_dpath_pmp_5_mask[20] : io_dpath_pmp_5_mask[29]; // @[package.scala 32:76]
  assign _T_756 = _T_44 ? io_dpath_pmp_5_mask[11] : _T_754; // @[package.scala 32:76]
  assign _T_758 = _T_46 ? io_dpath_pmp_5_mask[11] : _T_756; // @[package.scala 32:76]
  assign _T_759 = {io_dpath_pmp_5_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_761 = ~_T_759 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_159 = {{34'd0}, ~_T_761}; // @[PMP.scala 100:53]
  assign _T_763 = _T_357 ^ _GEN_159; // @[PMP.scala 100:53]
  assign _T_765 = _T_763[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _T_772 = _T_763[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _T_779 = _T_763[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _T_781 = _T_42 ? _T_772 : _T_765; // @[package.scala 32:76]
  assign _T_783 = _T_44 ? _T_779 : _T_781; // @[package.scala 32:76]
  assign _T_785 = _T_46 ? _T_779 : _T_783; // @[package.scala 32:76]
  assign _T_786 = _T_758 | _T_785; // @[PMP.scala 100:21]
  assign _T_799 = _T_357 < _GEN_159; // @[PMP.scala 109:32]
  assign _T_819 = ~_T_761 & _T_416; // @[PMP.scala 113:53]
  assign _GEN_167 = {{34'd0}, _T_819}; // @[PMP.scala 113:40]
  assign _T_820 = _T_417 < _GEN_167; // @[PMP.scala 113:40]
  assign _T_821 = _T_742 | ~_T_799; // @[PMP.scala 115:21]
  assign _T_822 = ~_T_721 & _T_820; // @[PMP.scala 115:62]
  assign _T_823 = _T_821 | _T_822; // @[PMP.scala 115:41]
  assign _T_824 = ~io_dpath_pmp_5_cfg_a[0] | _T_823; // @[PMP.scala 120:58]
  assign _T_825 = io_dpath_pmp_5_cfg_a[1] ? _T_786 : _T_824; // @[PMP.scala 120:8]
  assign _T_826 = _T_748 & _T_825; // @[PMP.scala 140:10]
  assign _T_832 = _T_42 ? io_dpath_pmp_6_mask[20] : io_dpath_pmp_6_mask[29]; // @[package.scala 32:76]
  assign _T_834 = _T_44 ? io_dpath_pmp_6_mask[11] : _T_832; // @[package.scala 32:76]
  assign _T_836 = _T_46 ? io_dpath_pmp_6_mask[11] : _T_834; // @[package.scala 32:76]
  assign _T_837 = {io_dpath_pmp_6_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_839 = ~_T_837 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_168 = {{34'd0}, ~_T_839}; // @[PMP.scala 100:53]
  assign _T_841 = _T_357 ^ _GEN_168; // @[PMP.scala 100:53]
  assign _T_843 = _T_841[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _T_850 = _T_841[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _T_857 = _T_841[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _T_859 = _T_42 ? _T_850 : _T_843; // @[package.scala 32:76]
  assign _T_861 = _T_44 ? _T_857 : _T_859; // @[package.scala 32:76]
  assign _T_863 = _T_46 ? _T_857 : _T_861; // @[package.scala 32:76]
  assign _T_864 = _T_836 | _T_863; // @[PMP.scala 100:21]
  assign _T_877 = _T_357 < _GEN_168; // @[PMP.scala 109:32]
  assign _T_897 = ~_T_839 & _T_416; // @[PMP.scala 113:53]
  assign _GEN_176 = {{34'd0}, _T_897}; // @[PMP.scala 113:40]
  assign _T_898 = _T_417 < _GEN_176; // @[PMP.scala 113:40]
  assign _T_899 = _T_820 | ~_T_877; // @[PMP.scala 115:21]
  assign _T_900 = ~_T_799 & _T_898; // @[PMP.scala 115:62]
  assign _T_901 = _T_899 | _T_900; // @[PMP.scala 115:41]
  assign _T_902 = ~io_dpath_pmp_6_cfg_a[0] | _T_901; // @[PMP.scala 120:58]
  assign _T_903 = io_dpath_pmp_6_cfg_a[1] ? _T_864 : _T_902; // @[PMP.scala 120:8]
  assign _T_904 = _T_826 & _T_903; // @[PMP.scala 140:10]
  assign _T_910 = _T_42 ? io_dpath_pmp_7_mask[20] : io_dpath_pmp_7_mask[29]; // @[package.scala 32:76]
  assign _T_912 = _T_44 ? io_dpath_pmp_7_mask[11] : _T_910; // @[package.scala 32:76]
  assign _T_914 = _T_46 ? io_dpath_pmp_7_mask[11] : _T_912; // @[package.scala 32:76]
  assign _T_915 = {io_dpath_pmp_7_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_917 = ~_T_915 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_177 = {{34'd0}, ~_T_917}; // @[PMP.scala 100:53]
  assign _T_919 = _T_357 ^ _GEN_177; // @[PMP.scala 100:53]
  assign _T_921 = _T_919[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _T_928 = _T_919[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _T_935 = _T_919[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _T_937 = _T_42 ? _T_928 : _T_921; // @[package.scala 32:76]
  assign _T_939 = _T_44 ? _T_935 : _T_937; // @[package.scala 32:76]
  assign _T_941 = _T_46 ? _T_935 : _T_939; // @[package.scala 32:76]
  assign _T_942 = _T_914 | _T_941; // @[PMP.scala 100:21]
  assign _T_955 = _T_357 < _GEN_177; // @[PMP.scala 109:32]
  assign _T_975 = ~_T_917 & _T_416; // @[PMP.scala 113:53]
  assign _GEN_185 = {{34'd0}, _T_975}; // @[PMP.scala 113:40]
  assign _T_976 = _T_417 < _GEN_185; // @[PMP.scala 113:40]
  assign _T_977 = _T_898 | ~_T_955; // @[PMP.scala 115:21]
  assign _T_978 = ~_T_877 & _T_976; // @[PMP.scala 115:62]
  assign _T_979 = _T_977 | _T_978; // @[PMP.scala 115:41]
  assign _T_980 = ~io_dpath_pmp_7_cfg_a[0] | _T_979; // @[PMP.scala 120:58]
  assign _T_981 = io_dpath_pmp_7_cfg_a[1] ? _T_942 : _T_980; // @[PMP.scala 120:8]
  assign pmpHomogeneous = _T_904 & _T_981; // @[PMP.scala 140:10]
  assign homogeneous = pmaHomogeneous & pmpHomogeneous; // @[PTW.scala 269:36]
  assign _T_986 = 3'h0 == state; // @[Conditional.scala 37:30]
  assign _T_988 = arb_io_out_bits_valid ? 3'h1 : 3'h0; // @[PTW.scala 291:26]
  assign _GEN_40 = _T_55 ? _T_988 : state; // @[PTW.scala 290:32]
  assign _T_990 = 1'h0 - 1'h0; // @[PTW.scala 293:39]
  assign _T_991 = 3'h1 == state; // @[Conditional.scala 37:30]
  assign _T_993 = count + 2'h1; // @[PTW.scala 297:24]
  assign _T_994 = io_mem_req_ready ? 3'h2 : 3'h1; // @[PTW.scala 299:26]
  assign _GEN_42 = pte_cache_hit ? state : _T_994; // @[PTW.scala 296:28]
  assign _T_995 = 3'h2 == state; // @[Conditional.scala 37:30]
  assign _T_997 = 3'h4 == state; // @[Conditional.scala 37:30]
  assign _GEN_46 = io_mem_s2_xcpt_ae_ld ? 3'h0 : 3'h5; // @[PTW.scala 308:35]
  assign _GEN_47 = io_mem_s2_xcpt_ae_ld & ~r_req_dest; // @[PTW.scala 308:35]
  assign _GEN_48 = io_mem_s2_xcpt_ae_ld & r_req_dest; // @[PTW.scala 308:35]
  assign _T_1000 = 3'h7 == state; // @[Conditional.scala 37:30]
  assign _GEN_53 = _T_1000 ? 3'h0 : state; // @[Conditional.scala 39:67]
  assign _GEN_54 = _T_1000 & ~r_req_dest; // @[Conditional.scala 39:67]
  assign _GEN_55 = _T_1000 & r_req_dest; // @[Conditional.scala 39:67]
  assign _GEN_59 = _T_997 ? _GEN_46 : _GEN_53; // @[Conditional.scala 39:67]
  assign _GEN_60 = _T_997 & io_mem_s2_xcpt_ae_ld; // @[Conditional.scala 39:67]
  assign _GEN_61 = _T_997 ? _GEN_47 : _GEN_54; // @[Conditional.scala 39:67]
  assign _GEN_62 = _T_997 ? _GEN_48 : _GEN_55; // @[Conditional.scala 39:67]
  assign _GEN_65 = _T_995 ? 3'h4 : _GEN_59; // @[Conditional.scala 39:67]
  assign _GEN_67 = _T_995 ? 1'h0 : _GEN_61; // @[Conditional.scala 39:67]
  assign _GEN_68 = _T_995 ? 1'h0 : _GEN_62; // @[Conditional.scala 39:67]
  assign _GEN_72 = _T_991 ? _GEN_42 : _GEN_65; // @[Conditional.scala 39:67]
  assign _GEN_74 = _T_991 ? 1'h0 : _GEN_67; // @[Conditional.scala 39:67]
  assign _GEN_75 = _T_991 ? 1'h0 : _GEN_68; // @[Conditional.scala 39:67]
  assign _GEN_77 = _T_986 ? _GEN_40 : _GEN_72; // @[Conditional.scala 40:58]
  assign _GEN_80 = _T_986 ? 1'h0 : _GEN_74; // @[Conditional.scala 40:58]
  assign _GEN_81 = _T_986 ? 1'h0 : _GEN_75; // @[Conditional.scala 40:58]
  assign _T_1006 = state == 3'h7; // @[PTW.scala 333:15]
  assign _T_1008 = _T_1006 & ~homogeneous; // @[PTW.scala 333:40]
  assign _T_1010 = _T_115 & pte_cache_hit; // @[PTW.scala 334:25]
  assign pte_2_ppn = {{10'd0}, io_dpath_ptbr_ppn}; // @[PTW.scala 327:13]
  assign _T_1012_ppn = _T_55 ? pte_2_ppn : r_pte_ppn; // @[PTW.scala 335:8]
  assign pte_1_ppn = {{34'd0}, pte_cache_data}; // @[PTW.scala 327:13]
  assign _T_1013_ppn = _T_1010 ? pte_1_ppn : _T_1012_ppn; // @[PTW.scala 334:8]
  assign _T_1013_d = _T_1010 ? 1'h0 : r_pte_d; // @[PTW.scala 334:8]
  assign _T_1013_a = _T_1010 ? 1'h0 : r_pte_a; // @[PTW.scala 334:8]
  assign _T_1013_g = _T_1010 ? 1'h0 : r_pte_g; // @[PTW.scala 334:8]
  assign _T_1013_u = _T_1010 ? 1'h0 : r_pte_u; // @[PTW.scala 334:8]
  assign _T_1013_x = _T_1010 ? 1'h0 : r_pte_x; // @[PTW.scala 334:8]
  assign _T_1013_w = _T_1010 ? 1'h0 : r_pte_w; // @[PTW.scala 334:8]
  assign _T_1013_r = _T_1010 ? 1'h0 : r_pte_r; // @[PTW.scala 334:8]
  assign _T_1013_v = _T_1010 ? 1'h0 : r_pte_v; // @[PTW.scala 334:8]
  assign _T_1014_ppn = _T_1008 ? fragmented_superpage_ppn : _T_1013_ppn; // @[PTW.scala 333:8]
  assign _T_1014_d = _T_1008 ? r_pte_d : _T_1013_d; // @[PTW.scala 333:8]
  assign _T_1014_a = _T_1008 ? r_pte_a : _T_1013_a; // @[PTW.scala 333:8]
  assign _T_1014_g = _T_1008 ? r_pte_g : _T_1013_g; // @[PTW.scala 333:8]
  assign _T_1014_u = _T_1008 ? r_pte_u : _T_1013_u; // @[PTW.scala 333:8]
  assign _T_1014_x = _T_1008 ? r_pte_x : _T_1013_x; // @[PTW.scala 333:8]
  assign _T_1014_w = _T_1008 ? r_pte_w : _T_1013_w; // @[PTW.scala 333:8]
  assign _T_1014_r = _T_1008 ? r_pte_r : _T_1013_r; // @[PTW.scala 333:8]
  assign _T_1014_v = _T_1008 ? r_pte_v : _T_1013_v; // @[PTW.scala 333:8]
  assign _GEN_83 = ~r_req_dest | _GEN_80; // @[PTW.scala 341:28]
  assign _GEN_84 = r_req_dest | _GEN_81; // @[PTW.scala 341:28]
  assign _T_1027 = state == 3'h5; // @[PTW.scala 346:18]
  assign _T_1029 = _T_1027 | reset; // @[PTW.scala 346:11]
  assign ae = res_v & invalid_paddr; // @[PTW.scala 352:22]
  assign _GEN_95 = traverse ? 3'h1 : 3'h0; // @[PTW.scala 347:21]
  assign _GEN_101 = mem_resp_valid ? _GEN_95 : _GEN_77; // @[PTW.scala 345:25]
  assign _T_1043 = state == 3'h4; // @[PTW.scala 363:18]
  assign _T_1045 = _T_1043 | reset; // @[PTW.scala 363:11]
  assign io_requestor_0_req_ready = arb_io_in_0_ready; // @[PTW.scala 106:13]
  assign io_requestor_0_resp_valid = resp_valid_0; // @[PTW.scala 272:32]
  assign io_requestor_0_resp_bits_ae = resp_ae; // @[PTW.scala 273:34]
  assign io_requestor_0_resp_bits_pte_ppn = r_pte_ppn; // @[PTW.scala 274:35]
  assign io_requestor_0_resp_bits_pte_d = r_pte_d; // @[PTW.scala 274:35]
  assign io_requestor_0_resp_bits_pte_a = r_pte_a; // @[PTW.scala 274:35]
  assign io_requestor_0_resp_bits_pte_g = r_pte_g; // @[PTW.scala 274:35]
  assign io_requestor_0_resp_bits_pte_u = r_pte_u; // @[PTW.scala 274:35]
  assign io_requestor_0_resp_bits_pte_x = r_pte_x; // @[PTW.scala 274:35]
  assign io_requestor_0_resp_bits_pte_w = r_pte_w; // @[PTW.scala 274:35]
  assign io_requestor_0_resp_bits_pte_r = r_pte_r; // @[PTW.scala 274:35]
  assign io_requestor_0_resp_bits_pte_v = r_pte_v; // @[PTW.scala 274:35]
  assign io_requestor_0_resp_bits_level = count; // @[PTW.scala 275:37]
  assign io_requestor_0_resp_bits_homogeneous = pmaHomogeneous & pmpHomogeneous; // @[PTW.scala 276:43]
  assign io_requestor_0_ptbr_mode = io_dpath_ptbr_mode; // @[PTW.scala 278:26]
  assign io_requestor_0_status_debug = io_dpath_status_debug; // @[PTW.scala 280:28]
  assign io_requestor_0_status_dprv = io_dpath_status_dprv; // @[PTW.scala 280:28]
  assign io_requestor_0_status_mxr = io_dpath_status_mxr; // @[PTW.scala 280:28]
  assign io_requestor_0_status_sum = io_dpath_status_sum; // @[PTW.scala 280:28]
  assign io_requestor_0_pmp_0_cfg_l = io_dpath_pmp_0_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_0_cfg_a = io_dpath_pmp_0_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_0_cfg_x = io_dpath_pmp_0_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_0_cfg_w = io_dpath_pmp_0_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_0_cfg_r = io_dpath_pmp_0_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_0_addr = io_dpath_pmp_0_addr; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_0_mask = io_dpath_pmp_0_mask; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_1_cfg_l = io_dpath_pmp_1_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_1_cfg_a = io_dpath_pmp_1_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_1_cfg_x = io_dpath_pmp_1_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_1_cfg_w = io_dpath_pmp_1_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_1_cfg_r = io_dpath_pmp_1_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_1_addr = io_dpath_pmp_1_addr; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_1_mask = io_dpath_pmp_1_mask; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_2_cfg_l = io_dpath_pmp_2_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_2_cfg_a = io_dpath_pmp_2_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_2_cfg_x = io_dpath_pmp_2_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_2_cfg_w = io_dpath_pmp_2_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_2_cfg_r = io_dpath_pmp_2_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_2_addr = io_dpath_pmp_2_addr; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_2_mask = io_dpath_pmp_2_mask; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_3_cfg_l = io_dpath_pmp_3_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_3_cfg_a = io_dpath_pmp_3_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_3_cfg_x = io_dpath_pmp_3_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_3_cfg_w = io_dpath_pmp_3_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_3_cfg_r = io_dpath_pmp_3_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_3_addr = io_dpath_pmp_3_addr; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_3_mask = io_dpath_pmp_3_mask; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_4_cfg_l = io_dpath_pmp_4_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_4_cfg_a = io_dpath_pmp_4_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_4_cfg_x = io_dpath_pmp_4_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_4_cfg_w = io_dpath_pmp_4_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_4_cfg_r = io_dpath_pmp_4_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_4_addr = io_dpath_pmp_4_addr; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_4_mask = io_dpath_pmp_4_mask; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_5_cfg_l = io_dpath_pmp_5_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_5_cfg_a = io_dpath_pmp_5_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_5_cfg_x = io_dpath_pmp_5_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_5_cfg_w = io_dpath_pmp_5_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_5_cfg_r = io_dpath_pmp_5_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_5_addr = io_dpath_pmp_5_addr; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_5_mask = io_dpath_pmp_5_mask; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_6_cfg_l = io_dpath_pmp_6_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_6_cfg_a = io_dpath_pmp_6_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_6_cfg_x = io_dpath_pmp_6_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_6_cfg_w = io_dpath_pmp_6_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_6_cfg_r = io_dpath_pmp_6_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_6_addr = io_dpath_pmp_6_addr; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_6_mask = io_dpath_pmp_6_mask; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_7_cfg_l = io_dpath_pmp_7_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_7_cfg_a = io_dpath_pmp_7_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_7_cfg_x = io_dpath_pmp_7_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_7_cfg_w = io_dpath_pmp_7_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_7_cfg_r = io_dpath_pmp_7_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_7_addr = io_dpath_pmp_7_addr; // @[PTW.scala 281:25]
  assign io_requestor_0_pmp_7_mask = io_dpath_pmp_7_mask; // @[PTW.scala 281:25]
  assign io_requestor_1_req_ready = arb_io_in_1_ready; // @[PTW.scala 106:13]
  assign io_requestor_1_resp_valid = resp_valid_1; // @[PTW.scala 272:32]
  assign io_requestor_1_resp_bits_ae = resp_ae; // @[PTW.scala 273:34]
  assign io_requestor_1_resp_bits_pte_ppn = r_pte_ppn; // @[PTW.scala 274:35]
  assign io_requestor_1_resp_bits_pte_d = r_pte_d; // @[PTW.scala 274:35]
  assign io_requestor_1_resp_bits_pte_a = r_pte_a; // @[PTW.scala 274:35]
  assign io_requestor_1_resp_bits_pte_g = r_pte_g; // @[PTW.scala 274:35]
  assign io_requestor_1_resp_bits_pte_u = r_pte_u; // @[PTW.scala 274:35]
  assign io_requestor_1_resp_bits_pte_x = r_pte_x; // @[PTW.scala 274:35]
  assign io_requestor_1_resp_bits_pte_w = r_pte_w; // @[PTW.scala 274:35]
  assign io_requestor_1_resp_bits_pte_r = r_pte_r; // @[PTW.scala 274:35]
  assign io_requestor_1_resp_bits_pte_v = r_pte_v; // @[PTW.scala 274:35]
  assign io_requestor_1_resp_bits_level = count; // @[PTW.scala 275:37]
  assign io_requestor_1_resp_bits_homogeneous = pmaHomogeneous & pmpHomogeneous; // @[PTW.scala 276:43]
  assign io_requestor_1_ptbr_mode = io_dpath_ptbr_mode; // @[PTW.scala 278:26]
  assign io_requestor_1_status_debug = io_dpath_status_debug; // @[PTW.scala 280:28]
  assign io_requestor_1_status_prv = io_dpath_status_prv; // @[PTW.scala 280:28]
  assign io_requestor_1_pmp_0_cfg_l = io_dpath_pmp_0_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_0_cfg_a = io_dpath_pmp_0_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_0_cfg_x = io_dpath_pmp_0_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_0_cfg_w = io_dpath_pmp_0_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_0_cfg_r = io_dpath_pmp_0_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_0_addr = io_dpath_pmp_0_addr; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_0_mask = io_dpath_pmp_0_mask; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_1_cfg_l = io_dpath_pmp_1_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_1_cfg_a = io_dpath_pmp_1_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_1_cfg_x = io_dpath_pmp_1_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_1_cfg_w = io_dpath_pmp_1_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_1_cfg_r = io_dpath_pmp_1_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_1_addr = io_dpath_pmp_1_addr; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_1_mask = io_dpath_pmp_1_mask; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_2_cfg_l = io_dpath_pmp_2_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_2_cfg_a = io_dpath_pmp_2_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_2_cfg_x = io_dpath_pmp_2_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_2_cfg_w = io_dpath_pmp_2_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_2_cfg_r = io_dpath_pmp_2_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_2_addr = io_dpath_pmp_2_addr; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_2_mask = io_dpath_pmp_2_mask; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_3_cfg_l = io_dpath_pmp_3_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_3_cfg_a = io_dpath_pmp_3_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_3_cfg_x = io_dpath_pmp_3_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_3_cfg_w = io_dpath_pmp_3_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_3_cfg_r = io_dpath_pmp_3_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_3_addr = io_dpath_pmp_3_addr; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_3_mask = io_dpath_pmp_3_mask; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_4_cfg_l = io_dpath_pmp_4_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_4_cfg_a = io_dpath_pmp_4_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_4_cfg_x = io_dpath_pmp_4_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_4_cfg_w = io_dpath_pmp_4_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_4_cfg_r = io_dpath_pmp_4_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_4_addr = io_dpath_pmp_4_addr; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_4_mask = io_dpath_pmp_4_mask; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_5_cfg_l = io_dpath_pmp_5_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_5_cfg_a = io_dpath_pmp_5_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_5_cfg_x = io_dpath_pmp_5_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_5_cfg_w = io_dpath_pmp_5_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_5_cfg_r = io_dpath_pmp_5_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_5_addr = io_dpath_pmp_5_addr; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_5_mask = io_dpath_pmp_5_mask; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_6_cfg_l = io_dpath_pmp_6_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_6_cfg_a = io_dpath_pmp_6_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_6_cfg_x = io_dpath_pmp_6_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_6_cfg_w = io_dpath_pmp_6_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_6_cfg_r = io_dpath_pmp_6_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_6_addr = io_dpath_pmp_6_addr; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_6_mask = io_dpath_pmp_6_mask; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_7_cfg_l = io_dpath_pmp_7_cfg_l; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_7_cfg_a = io_dpath_pmp_7_cfg_a; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_7_cfg_x = io_dpath_pmp_7_cfg_x; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_7_cfg_w = io_dpath_pmp_7_cfg_w; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_7_cfg_r = io_dpath_pmp_7_cfg_r; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_7_addr = io_dpath_pmp_7_addr; // @[PTW.scala 281:25]
  assign io_requestor_1_pmp_7_mask = io_dpath_pmp_7_mask; // @[PTW.scala 281:25]
  assign io_requestor_1_customCSRs_csrs_0_value = io_dpath_customCSRs_csrs_0_value; // @[PTW.scala 279:32]
  assign io_mem_req_valid = _T_115 | _T_205; // @[PTW.scala 247:20]
  assign io_mem_req_bits_addr = pte_addr[39:0]; // @[PTW.scala 252:24]
  assign io_mem_s1_kill = state != 3'h2; // @[PTW.scala 254:18]
  assign arb_io_in_0_valid = io_requestor_0_req_valid; // @[PTW.scala 106:13]
  assign arb_io_in_0_bits_bits_addr = io_requestor_0_req_bits_bits_addr; // @[PTW.scala 106:13]
  assign arb_io_in_1_valid = io_requestor_1_req_valid; // @[PTW.scala 106:13]
  assign arb_io_in_1_bits_valid = io_requestor_1_req_bits_valid; // @[PTW.scala 106:13]
  assign arb_io_in_1_bits_bits_addr = io_requestor_1_req_bits_bits_addr; // @[PTW.scala 106:13]
  assign arb_io_out_ready = state == 3'h0; // @[PTW.scala 107:20]
  assign OptimizationBarrier_io_x = io_mem_s2_nack ? 3'h1 : _GEN_101; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_ppn = mem_resp_valid ? res_ppn : _T_1014_ppn; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_d = mem_resp_valid ? tmp_d : _T_1014_d; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_a = mem_resp_valid ? tmp_a : _T_1014_a; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_g = mem_resp_valid ? tmp_g : _T_1014_g; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_u = mem_resp_valid ? tmp_u : _T_1014_u; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_x = mem_resp_valid ? tmp_x : _T_1014_x; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_w = mem_resp_valid ? tmp_w : _T_1014_w; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_r = mem_resp_valid ? tmp_r : _T_1014_r; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_v = mem_resp_valid ? res_v : _T_1014_v; // @[package.scala 244:18]
  assign PTW_cov_read_addr = PTW_state;
  assign PTW_cov_read_data = PTW_cov[PTW_cov_read_addr]; // @[Coverage map for PTW]
  assign PTW_cov_write_data = 1'h1;
  assign PTW_cov_write_addr = PTW_state;
  assign PTW_cov_write_mask = 1'h1;
  assign PTW_cov_write_en = 1'h1;
  assign valid_shl = {valid, 3'h0};
  assign valid_pad = {9'h0,valid_shl};
  assign invalidated_shl = {invalidated, 11'h0};
  assign invalidated_pad = {8'h0,invalidated_shl};
  assign state_shl = {state, 10'h0};
  assign state_pad = {7'h0,state_shl};
  assign _T_56_shl = _T_56;
  assign _T_56_pad = {13'h0,_T_56_shl};
  assign count_shl = {count, 14'h0};
  assign count_pad = {4'h0,count_shl};
  assign mem_resp_valid_shl = {mem_resp_valid, 1'h0};
  assign mem_resp_valid_pad = {18'h0,mem_resp_valid_shl};
  assign PTW_xor4 = invalidated_pad ^ state_pad;
  assign PTW_xor1 = valid_pad ^ PTW_xor4;
  assign PTW_xor6 = count_pad ^ mem_resp_valid_pad;
  assign PTW_xor2 = _T_56_pad ^ PTW_xor6;
  assign PTW_xor0 = PTW_xor1 ^ PTW_xor2;
  assign arb_sum = PTW_covSum + arb_io_covSum;
  assign OptimizationBarrier_sum = arb_sum + OptimizationBarrier_io_covSum;
  assign OptimizationBarrier_1_sum = OptimizationBarrier_sum + OptimizationBarrier_1_io_covSum;
  assign io_covSum = OptimizationBarrier_1_sum;
  assign stopEn0 = mem_resp_valid & ~_T_1029;
  assign stopEn1 = io_mem_s2_nack & ~_T_1045;
  assign arb_metaAssert_wire = arb_metaAssert;
  assign OptimizationBarrier_metaAssert_wire = OptimizationBarrier_metaAssert;
  assign OptimizationBarrier_1_metaAssert_wire = OptimizationBarrier_1_metaAssert;
  assign PTW_or1 = stopEn0 | stopEn1;
  assign PTW_or6 = OptimizationBarrier_metaAssert_wire | OptimizationBarrier_1_metaAssert_wire;
  assign PTW_or2 = arb_metaAssert_wire | PTW_or6;
  assign PTW_or0 = PTW_or1 | PTW_or2;
  assign metaAssert = PTW_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  resp_valid_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  resp_valid_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  invalidated = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  count = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  resp_ae = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  r_req_addr = _RAND_6[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  r_req_dest = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  r_pte_ppn = _RAND_8[53:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  r_pte_d = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  r_pte_a = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  r_pte_g = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  r_pte_u = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  r_pte_x = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  r_pte_w = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  r_pte_r = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  r_pte_v = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  mem_resp_valid = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  mem_resp_data = _RAND_18[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_56 = _RAND_19[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  valid = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  tags_0 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  tags_1 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  tags_2 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  tags_3 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  tags_4 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  tags_5 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  tags_6 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  tags_7 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  data_0 = _RAND_29[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  data_1 = _RAND_30[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  data_2 = _RAND_31[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  data_3 = _RAND_32[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  data_4 = _RAND_33[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  data_5 = _RAND_34[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  data_6 = _RAND_35[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  data_7 = _RAND_36[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  PTW_state = _RAND_37[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    PTW_cov[initvar] = _RAND_38[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  PTW_covSum = _RAND_39[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  PTW_metaAssert = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      state <= 3'h0;
    end else if (reset) begin
      state <= 3'h0;
    end else begin
      state <= OptimizationBarrier_io_y;
    end
    if (metaReset) begin
      resp_valid_0 <= 1'h0;
    end else if (mem_resp_valid) begin
      if (traverse) begin
        if (_T_986) begin
          resp_valid_0 <= 1'h0;
        end else if (_T_991) begin
          resp_valid_0 <= 1'h0;
        end else if (_T_995) begin
          resp_valid_0 <= 1'h0;
        end else if (_T_997) begin
          resp_valid_0 <= _GEN_47;
        end else begin
          resp_valid_0 <= _GEN_54;
        end
      end else begin
        resp_valid_0 <= _GEN_83;
      end
    end else if (_T_986) begin
      resp_valid_0 <= 1'h0;
    end else if (_T_991) begin
      resp_valid_0 <= 1'h0;
    end else if (_T_995) begin
      resp_valid_0 <= 1'h0;
    end else if (_T_997) begin
      resp_valid_0 <= _GEN_47;
    end else begin
      resp_valid_0 <= _GEN_54;
    end
    if (metaReset) begin
      resp_valid_1 <= 1'h0;
    end else if (mem_resp_valid) begin
      if (traverse) begin
        if (_T_986) begin
          resp_valid_1 <= 1'h0;
        end else if (_T_991) begin
          resp_valid_1 <= 1'h0;
        end else if (_T_995) begin
          resp_valid_1 <= 1'h0;
        end else if (_T_997) begin
          resp_valid_1 <= _GEN_48;
        end else begin
          resp_valid_1 <= _GEN_55;
        end
      end else begin
        resp_valid_1 <= _GEN_84;
      end
    end else if (_T_986) begin
      resp_valid_1 <= 1'h0;
    end else if (_T_991) begin
      resp_valid_1 <= 1'h0;
    end else if (_T_995) begin
      resp_valid_1 <= 1'h0;
    end else if (_T_997) begin
      resp_valid_1 <= _GEN_48;
    end else begin
      resp_valid_1 <= _GEN_55;
    end
    if (metaReset) begin
      invalidated <= 1'h0;
    end else begin
      invalidated <= io_dpath_sfence_valid | _T_202;
    end
    if (metaReset) begin
      count <= 2'h0;
    end else if (mem_resp_valid) begin
      if (traverse) begin
        count <= _T_993;
      end else if (_T_986) begin
        count <= {{1'd0}, _T_990};
      end else if (_T_991) begin
        if (pte_cache_hit) begin
          count <= _T_993;
        end
      end else if (!(_T_995)) begin
        if (!(_T_997)) begin
          if (_T_1000) begin
            if (~homogeneous) begin
              count <= 2'h2;
            end
          end
        end
      end
    end else if (_T_986) begin
      count <= {{1'd0}, _T_990};
    end else if (_T_991) begin
      if (pte_cache_hit) begin
        count <= _T_993;
      end
    end else if (!(_T_995)) begin
      if (!(_T_997)) begin
        if (_T_1000) begin
          if (~homogeneous) begin
            count <= 2'h2;
          end
        end
      end
    end
    if (metaReset) begin
      resp_ae <= 1'h0;
    end else if (mem_resp_valid) begin
      if (traverse) begin
        if (_T_986) begin
          resp_ae <= 1'h0;
        end else if (_T_991) begin
          resp_ae <= 1'h0;
        end else if (_T_995) begin
          resp_ae <= 1'h0;
        end else begin
          resp_ae <= _GEN_60;
        end
      end else begin
        resp_ae <= ae;
      end
    end else if (_T_986) begin
      resp_ae <= 1'h0;
    end else if (_T_991) begin
      resp_ae <= 1'h0;
    end else if (_T_995) begin
      resp_ae <= 1'h0;
    end else begin
      resp_ae <= _GEN_60;
    end
    if (metaReset) begin
      r_req_addr <= 27'h0;
    end else if (_T_55) begin
      r_req_addr <= arb_io_out_bits_bits_addr;
    end
    if (metaReset) begin
      r_req_dest <= 1'h0;
    end else if (_T_55) begin
      r_req_dest <= arb_io_chosen;
    end
    if (metaReset) begin
      r_pte_ppn <= 54'h0;
    end else begin
      r_pte_ppn <= OptimizationBarrier_1_io_y_ppn;
    end
    if (metaReset) begin
      r_pte_d <= 1'h0;
    end else begin
      r_pte_d <= OptimizationBarrier_1_io_y_d;
    end
    if (metaReset) begin
      r_pte_a <= 1'h0;
    end else begin
      r_pte_a <= OptimizationBarrier_1_io_y_a;
    end
    if (metaReset) begin
      r_pte_g <= 1'h0;
    end else begin
      r_pte_g <= OptimizationBarrier_1_io_y_g;
    end
    if (metaReset) begin
      r_pte_u <= 1'h0;
    end else begin
      r_pte_u <= OptimizationBarrier_1_io_y_u;
    end
    if (metaReset) begin
      r_pte_x <= 1'h0;
    end else begin
      r_pte_x <= OptimizationBarrier_1_io_y_x;
    end
    if (metaReset) begin
      r_pte_w <= 1'h0;
    end else begin
      r_pte_w <= OptimizationBarrier_1_io_y_w;
    end
    if (metaReset) begin
      r_pte_r <= 1'h0;
    end else begin
      r_pte_r <= OptimizationBarrier_1_io_y_r;
    end
    if (metaReset) begin
      r_pte_v <= 1'h0;
    end else begin
      r_pte_v <= OptimizationBarrier_1_io_y_v;
    end
    if (metaReset) begin
      mem_resp_valid <= 1'h0;
    end else begin
      mem_resp_valid <= io_mem_resp_valid;
    end
    if (metaReset) begin
      mem_resp_data <= 64'h0;
    end else begin
      mem_resp_data <= io_mem_resp_bits_data;
    end
    if (metaReset) begin
      _T_56 <= 7'h0;
    end else if (_T_116) begin
      _T_56 <= _T_166;
    end
    if (metaReset) begin
      valid <= 8'h0;
    end else if (reset) begin
      valid <= 8'h0;
    end else if (_T_168) begin
      valid <= 8'h0;
    end else if (_T_76) begin
      valid <= _T_114;
    end
    if (metaReset) begin
      tags_0 <= 32'h0;
    end else if (_T_76) begin
      if (3'h0 == r) begin
        tags_0 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_1 <= 32'h0;
    end else if (_T_76) begin
      if (3'h1 == r) begin
        tags_1 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_2 <= 32'h0;
    end else if (_T_76) begin
      if (3'h2 == r) begin
        tags_2 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_3 <= 32'h0;
    end else if (_T_76) begin
      if (3'h3 == r) begin
        tags_3 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_4 <= 32'h0;
    end else if (_T_76) begin
      if (3'h4 == r) begin
        tags_4 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_5 <= 32'h0;
    end else if (_T_76) begin
      if (3'h5 == r) begin
        tags_5 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_6 <= 32'h0;
    end else if (_T_76) begin
      if (3'h6 == r) begin
        tags_6 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_7 <= 32'h0;
    end else if (_T_76) begin
      if (3'h7 == r) begin
        tags_7 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      data_0 <= 20'h0;
    end else if (_T_76) begin
      if (3'h0 == r) begin
        data_0 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_1 <= 20'h0;
    end else if (_T_76) begin
      if (3'h1 == r) begin
        data_1 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_2 <= 20'h0;
    end else if (_T_76) begin
      if (3'h2 == r) begin
        data_2 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_3 <= 20'h0;
    end else if (_T_76) begin
      if (3'h3 == r) begin
        data_3 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_4 <= 20'h0;
    end else if (_T_76) begin
      if (3'h4 == r) begin
        data_4 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_5 <= 20'h0;
    end else if (_T_76) begin
      if (3'h5 == r) begin
        data_5 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_6 <= 20'h0;
    end else if (_T_76) begin
      if (3'h6 == r) begin
        data_6 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_7 <= 20'h0;
    end else if (_T_76) begin
      if (3'h7 == r) begin
        data_7 <= res_ppn[19:0];
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (mem_resp_valid & ~_T_1029) begin
          $fwrite(32'h80000002,"Assertion failed\n    at PTW.scala:346 assert(state === s_wait3)\n"); // @[PTW.scala 346:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (mem_resp_valid & ~_T_1029) begin
          $fatal; // @[PTW.scala 346:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_mem_s2_nack & ~_T_1045) begin
          $fwrite(32'h80000002,"Assertion failed\n    at PTW.scala:363 assert(state === s_wait2)\n"); // @[PTW.scala 363:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_mem_s2_nack & ~_T_1045) begin
          $fatal; // @[PTW.scala 363:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    PTW_state <= PTW_xor0;
    if (!(PTW_cov_read_data)) begin
      PTW_covSum <= PTW_covSum + 1'h1;
    end
    if (metaReset) begin
      PTW_metaAssert <= 1'h0;
    end else begin
      PTW_metaAssert <= PTW_metaAssert | PTW_or0;
    end
  end
  always @(posedge clock) begin
    if(PTW_cov_write_en & PTW_cov_write_mask) begin
      PTW_cov[PTW_cov_write_addr] <= PTW_cov_write_data; // @[Coverage map for PTW]
    end
  end
endmodule
module Rocket(
  input         clock,
  input         reset,
  input         io_hartid,
  input         io_interrupts_debug,
  input         io_interrupts_mtip,
  input         io_interrupts_msip,
  input         io_interrupts_meip,
  input         io_interrupts_seip,
  output        io_imem_might_request,
  output        io_imem_req_valid,
  output [39:0] io_imem_req_bits_pc,
  output        io_imem_req_bits_speculative,
  output        io_imem_sfence_valid,
  output        io_imem_sfence_bits_rs1,
  output        io_imem_sfence_bits_rs2,
  output [38:0] io_imem_sfence_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input         io_imem_resp_bits_btb_taken,
  input         io_imem_resp_bits_btb_bridx,
  input  [4:0]  io_imem_resp_bits_btb_entry,
  input  [7:0]  io_imem_resp_bits_btb_bht_history,
  input  [39:0] io_imem_resp_bits_pc,
  input  [31:0] io_imem_resp_bits_data,
  input         io_imem_resp_bits_xcpt_pf_inst,
  input         io_imem_resp_bits_xcpt_ae_inst,
  input         io_imem_resp_bits_replay,
  output        io_imem_btb_update_valid,
  output [4:0]  io_imem_btb_update_bits_prediction_entry,
  output [38:0] io_imem_btb_update_bits_pc,
  output        io_imem_btb_update_bits_isValid,
  output [38:0] io_imem_btb_update_bits_br_pc,
  output [1:0]  io_imem_btb_update_bits_cfiType,
  output        io_imem_bht_update_valid,
  output [7:0]  io_imem_bht_update_bits_prediction_history,
  output [38:0] io_imem_bht_update_bits_pc,
  output        io_imem_bht_update_bits_branch,
  output        io_imem_bht_update_bits_taken,
  output        io_imem_bht_update_bits_mispredict,
  output        io_imem_flush_icache,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [39:0] io_dmem_req_bits_addr,
  output [6:0]  io_dmem_req_bits_tag,
  output [4:0]  io_dmem_req_bits_cmd,
  output [1:0]  io_dmem_req_bits_size,
  output        io_dmem_req_bits_signed,
  output        io_dmem_s1_kill,
  output [63:0] io_dmem_s1_data_data,
  input         io_dmem_s2_nack,
  input         io_dmem_resp_valid,
  input  [6:0]  io_dmem_resp_bits_tag,
  input  [1:0]  io_dmem_resp_bits_size,
  input  [63:0] io_dmem_resp_bits_data,
  input         io_dmem_resp_bits_replay,
  input         io_dmem_resp_bits_has_data,
  input  [63:0] io_dmem_resp_bits_data_word_bypass,
  input         io_dmem_replay_next,
  input         io_dmem_s2_xcpt_ma_ld,
  input         io_dmem_s2_xcpt_ma_st,
  input         io_dmem_s2_xcpt_pf_ld,
  input         io_dmem_s2_xcpt_pf_st,
  input         io_dmem_s2_xcpt_ae_ld,
  input         io_dmem_s2_xcpt_ae_st,
  input         io_dmem_ordered,
  input         io_dmem_perf_release,
  input         io_dmem_perf_grant,
  output [3:0]  io_ptw_ptbr_mode,
  output [43:0] io_ptw_ptbr_ppn,
  output        io_ptw_sfence_valid,
  output        io_ptw_sfence_bits_rs1,
  output        io_ptw_status_debug,
  output [1:0]  io_ptw_status_dprv,
  output [1:0]  io_ptw_status_prv,
  output        io_ptw_status_mxr,
  output        io_ptw_status_sum,
  output        io_ptw_pmp_0_cfg_l,
  output [1:0]  io_ptw_pmp_0_cfg_a,
  output        io_ptw_pmp_0_cfg_x,
  output        io_ptw_pmp_0_cfg_w,
  output        io_ptw_pmp_0_cfg_r,
  output [29:0] io_ptw_pmp_0_addr,
  output [31:0] io_ptw_pmp_0_mask,
  output        io_ptw_pmp_1_cfg_l,
  output [1:0]  io_ptw_pmp_1_cfg_a,
  output        io_ptw_pmp_1_cfg_x,
  output        io_ptw_pmp_1_cfg_w,
  output        io_ptw_pmp_1_cfg_r,
  output [29:0] io_ptw_pmp_1_addr,
  output [31:0] io_ptw_pmp_1_mask,
  output        io_ptw_pmp_2_cfg_l,
  output [1:0]  io_ptw_pmp_2_cfg_a,
  output        io_ptw_pmp_2_cfg_x,
  output        io_ptw_pmp_2_cfg_w,
  output        io_ptw_pmp_2_cfg_r,
  output [29:0] io_ptw_pmp_2_addr,
  output [31:0] io_ptw_pmp_2_mask,
  output        io_ptw_pmp_3_cfg_l,
  output [1:0]  io_ptw_pmp_3_cfg_a,
  output        io_ptw_pmp_3_cfg_x,
  output        io_ptw_pmp_3_cfg_w,
  output        io_ptw_pmp_3_cfg_r,
  output [29:0] io_ptw_pmp_3_addr,
  output [31:0] io_ptw_pmp_3_mask,
  output        io_ptw_pmp_4_cfg_l,
  output [1:0]  io_ptw_pmp_4_cfg_a,
  output        io_ptw_pmp_4_cfg_x,
  output        io_ptw_pmp_4_cfg_w,
  output        io_ptw_pmp_4_cfg_r,
  output [29:0] io_ptw_pmp_4_addr,
  output [31:0] io_ptw_pmp_4_mask,
  output        io_ptw_pmp_5_cfg_l,
  output [1:0]  io_ptw_pmp_5_cfg_a,
  output        io_ptw_pmp_5_cfg_x,
  output        io_ptw_pmp_5_cfg_w,
  output        io_ptw_pmp_5_cfg_r,
  output [29:0] io_ptw_pmp_5_addr,
  output [31:0] io_ptw_pmp_5_mask,
  output        io_ptw_pmp_6_cfg_l,
  output [1:0]  io_ptw_pmp_6_cfg_a,
  output        io_ptw_pmp_6_cfg_x,
  output        io_ptw_pmp_6_cfg_w,
  output        io_ptw_pmp_6_cfg_r,
  output [29:0] io_ptw_pmp_6_addr,
  output [31:0] io_ptw_pmp_6_mask,
  output        io_ptw_pmp_7_cfg_l,
  output [1:0]  io_ptw_pmp_7_cfg_a,
  output        io_ptw_pmp_7_cfg_x,
  output        io_ptw_pmp_7_cfg_w,
  output        io_ptw_pmp_7_cfg_r,
  output [29:0] io_ptw_pmp_7_addr,
  output [31:0] io_ptw_pmp_7_mask,
  output [63:0] io_ptw_customCSRs_csrs_0_value,
  output [31:0] io_fpu_inst,
  output [63:0] io_fpu_fromint_data,
  output [2:0]  io_fpu_fcsr_rm,
  input         io_fpu_fcsr_flags_valid,
  input  [4:0]  io_fpu_fcsr_flags_bits,
  input  [63:0] io_fpu_store_data,
  input  [63:0] io_fpu_toint_data,
  output        io_fpu_dmem_resp_val,
  output [2:0]  io_fpu_dmem_resp_type,
  output [4:0]  io_fpu_dmem_resp_tag,
  output [63:0] io_fpu_dmem_resp_data,
  output        io_fpu_valid,
  input         io_fpu_fcsr_rdy,
  input         io_fpu_nack_mem,
  input         io_fpu_illegal_rm,
  output        io_fpu_killx,
  output        io_fpu_killm,
  input         io_fpu_dec_wen,
  input         io_fpu_dec_ren1,
  input         io_fpu_dec_ren2,
  input         io_fpu_dec_ren3,
  input         io_fpu_sboard_set,
  input         io_fpu_sboard_clr,
  input  [4:0]  io_fpu_sboard_clra,
  output        io_wfi,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         csr_halt,
  input         div_halt,
  input         ibuf_halt,
  output [19:0] Checking_Rocket_regstate,	//Jaewon_Rocket_regstate
  output [29:0] Checking_Rocket_covSum	//Jaewon_Rocket_regstate
);
  assign Checking_Rocket_regstate = Rocket_state; 	//Jaewon_Rocket_regstate
  assign Checking_Rocket_covSum = Rocket_covSum; 	//Jaewon_Rocket_regstate
  wire  ibuf_clock; // @[RocketCore.scala 248:20]
  wire  ibuf_reset; // @[RocketCore.scala 248:20]
  wire  ibuf_io_imem_ready; // @[RocketCore.scala 248:20]
  wire  ibuf_io_imem_valid; // @[RocketCore.scala 248:20]
  wire  ibuf_io_imem_bits_btb_taken; // @[RocketCore.scala 248:20]
  wire  ibuf_io_imem_bits_btb_bridx; // @[RocketCore.scala 248:20]
  wire [4:0] ibuf_io_imem_bits_btb_entry; // @[RocketCore.scala 248:20]
  wire [7:0] ibuf_io_imem_bits_btb_bht_history; // @[RocketCore.scala 248:20]
  wire [39:0] ibuf_io_imem_bits_pc; // @[RocketCore.scala 248:20]
  wire [31:0] ibuf_io_imem_bits_data; // @[RocketCore.scala 248:20]
  wire  ibuf_io_imem_bits_xcpt_pf_inst; // @[RocketCore.scala 248:20]
  wire  ibuf_io_imem_bits_xcpt_ae_inst; // @[RocketCore.scala 248:20]
  wire  ibuf_io_imem_bits_replay; // @[RocketCore.scala 248:20]
  wire  ibuf_io_kill; // @[RocketCore.scala 248:20]
  wire [39:0] ibuf_io_pc; // @[RocketCore.scala 248:20]
  wire [4:0] ibuf_io_btb_resp_entry; // @[RocketCore.scala 248:20]
  wire [7:0] ibuf_io_btb_resp_bht_history; // @[RocketCore.scala 248:20]
  wire  ibuf_io_inst_0_ready; // @[RocketCore.scala 248:20]
  wire  ibuf_io_inst_0_valid; // @[RocketCore.scala 248:20]
  wire  ibuf_io_inst_0_bits_xcpt0_pf_inst; // @[RocketCore.scala 248:20]
  wire  ibuf_io_inst_0_bits_xcpt0_ae_inst; // @[RocketCore.scala 248:20]
  wire  ibuf_io_inst_0_bits_xcpt1_pf_inst; // @[RocketCore.scala 248:20]
  wire  ibuf_io_inst_0_bits_xcpt1_ae_inst; // @[RocketCore.scala 248:20]
  wire  ibuf_io_inst_0_bits_replay; // @[RocketCore.scala 248:20]
  wire  ibuf_io_inst_0_bits_rvc; // @[RocketCore.scala 248:20]
  wire [31:0] ibuf_io_inst_0_bits_inst_bits; // @[RocketCore.scala 248:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rd; // @[RocketCore.scala 248:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 248:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 248:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rs3; // @[RocketCore.scala 248:20]
  wire [31:0] ibuf_io_inst_0_bits_raw; // @[RocketCore.scala 248:20]
  wire [29:0] ibuf_io_covSum; // @[RocketCore.scala 248:20]
  wire  ibuf_metaAssert; // @[RocketCore.scala 248:20]
  wire  ibuf_metaReset; // @[RocketCore.scala 248:20]
  reg [63:0] _T_815 [0:30]; // @[RocketCore.scala 1014:15]
  reg [63:0] _RAND_0;
  wire [63:0] _T_815__T_820_data; // @[RocketCore.scala 1014:15]
  wire [4:0] _T_815__T_820_addr; // @[RocketCore.scala 1014:15]
  reg [63:0] _RAND_1;
  wire [63:0] _T_815__T_826_data; // @[RocketCore.scala 1014:15]
  wire [4:0] _T_815__T_826_addr; // @[RocketCore.scala 1014:15]
  reg [63:0] _RAND_2;
  wire [63:0] _T_815__T_1524_data; // @[RocketCore.scala 1014:15]
  wire [4:0] _T_815__T_1524_addr; // @[RocketCore.scala 1014:15]
  wire  _T_815__T_1524_mask; // @[RocketCore.scala 1014:15]
  wire  _T_815__T_1524_en; // @[RocketCore.scala 1014:15]
  wire  csr_clock; // @[RocketCore.scala 276:19]
  wire  csr_reset; // @[RocketCore.scala 276:19]
  wire  csr_io_ungated_clock; // @[RocketCore.scala 276:19]
  wire  csr_io_interrupts_debug; // @[RocketCore.scala 276:19]
  wire  csr_io_interrupts_mtip; // @[RocketCore.scala 276:19]
  wire  csr_io_interrupts_msip; // @[RocketCore.scala 276:19]
  wire  csr_io_interrupts_meip; // @[RocketCore.scala 276:19]
  wire  csr_io_interrupts_seip; // @[RocketCore.scala 276:19]
  wire  csr_io_hartid; // @[RocketCore.scala 276:19]
  wire [11:0] csr_io_rw_addr; // @[RocketCore.scala 276:19]
  wire [2:0] csr_io_rw_cmd; // @[RocketCore.scala 276:19]
  wire [63:0] csr_io_rw_rdata; // @[RocketCore.scala 276:19]
  wire [63:0] csr_io_rw_wdata; // @[RocketCore.scala 276:19]
  wire [11:0] csr_io_decode_0_csr; // @[RocketCore.scala 276:19]
  wire  csr_io_decode_0_fp_illegal; // @[RocketCore.scala 276:19]
  wire  csr_io_decode_0_fp_csr; // @[RocketCore.scala 276:19]
  wire  csr_io_decode_0_read_illegal; // @[RocketCore.scala 276:19]
  wire  csr_io_decode_0_write_illegal; // @[RocketCore.scala 276:19]
  wire  csr_io_decode_0_write_flush; // @[RocketCore.scala 276:19]
  wire  csr_io_decode_0_system_illegal; // @[RocketCore.scala 276:19]
  wire  csr_io_csr_stall; // @[RocketCore.scala 276:19]
  wire  csr_io_eret; // @[RocketCore.scala 276:19]
  wire  csr_io_singleStep; // @[RocketCore.scala 276:19]
  wire  csr_io_status_debug; // @[RocketCore.scala 276:19]
  wire  csr_io_status_cease; // @[RocketCore.scala 276:19]
  wire  csr_io_status_wfi; // @[RocketCore.scala 276:19]
  wire [31:0] csr_io_status_isa; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_status_dprv; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_status_prv; // @[RocketCore.scala 276:19]
  wire  csr_io_status_sd; // @[RocketCore.scala 276:19]
  wire [26:0] csr_io_status_zero2; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_status_sxl; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_status_uxl; // @[RocketCore.scala 276:19]
  wire  csr_io_status_sd_rv32; // @[RocketCore.scala 276:19]
  wire [7:0] csr_io_status_zero1; // @[RocketCore.scala 276:19]
  wire  csr_io_status_tsr; // @[RocketCore.scala 276:19]
  wire  csr_io_status_tw; // @[RocketCore.scala 276:19]
  wire  csr_io_status_tvm; // @[RocketCore.scala 276:19]
  wire  csr_io_status_mxr; // @[RocketCore.scala 276:19]
  wire  csr_io_status_sum; // @[RocketCore.scala 276:19]
  wire  csr_io_status_mprv; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_status_xs; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_status_fs; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_status_mpp; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_status_vs; // @[RocketCore.scala 276:19]
  wire  csr_io_status_spp; // @[RocketCore.scala 276:19]
  wire  csr_io_status_mpie; // @[RocketCore.scala 276:19]
  wire  csr_io_status_hpie; // @[RocketCore.scala 276:19]
  wire  csr_io_status_spie; // @[RocketCore.scala 276:19]
  wire  csr_io_status_upie; // @[RocketCore.scala 276:19]
  wire  csr_io_status_mie; // @[RocketCore.scala 276:19]
  wire  csr_io_status_hie; // @[RocketCore.scala 276:19]
  wire  csr_io_status_sie; // @[RocketCore.scala 276:19]
  wire  csr_io_status_uie; // @[RocketCore.scala 276:19]
  wire [3:0] csr_io_ptbr_mode; // @[RocketCore.scala 276:19]
  wire [43:0] csr_io_ptbr_ppn; // @[RocketCore.scala 276:19]
  wire [39:0] csr_io_evec; // @[RocketCore.scala 276:19]
  wire  csr_io_exception; // @[RocketCore.scala 276:19]
  wire  csr_io_retire; // @[RocketCore.scala 276:19]
  wire [63:0] csr_io_cause; // @[RocketCore.scala 276:19]
  wire [39:0] csr_io_pc; // @[RocketCore.scala 276:19]
  wire [39:0] csr_io_tval; // @[RocketCore.scala 276:19]
  wire [63:0] csr_io_time; // @[RocketCore.scala 276:19]
  wire [2:0] csr_io_fcsr_rm; // @[RocketCore.scala 276:19]
  wire  csr_io_fcsr_flags_valid; // @[RocketCore.scala 276:19]
  wire [4:0] csr_io_fcsr_flags_bits; // @[RocketCore.scala 276:19]
  wire  csr_io_interrupt; // @[RocketCore.scala 276:19]
  wire [63:0] csr_io_interrupt_cause; // @[RocketCore.scala 276:19]
  wire  csr_io_bp_0_control_action; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_bp_0_control_tmatch; // @[RocketCore.scala 276:19]
  wire  csr_io_bp_0_control_m; // @[RocketCore.scala 276:19]
  wire  csr_io_bp_0_control_s; // @[RocketCore.scala 276:19]
  wire  csr_io_bp_0_control_u; // @[RocketCore.scala 276:19]
  wire  csr_io_bp_0_control_x; // @[RocketCore.scala 276:19]
  wire  csr_io_bp_0_control_w; // @[RocketCore.scala 276:19]
  wire  csr_io_bp_0_control_r; // @[RocketCore.scala 276:19]
  wire [38:0] csr_io_bp_0_address; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_0_cfg_l; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_pmp_0_cfg_a; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_0_cfg_x; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_0_cfg_w; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_0_cfg_r; // @[RocketCore.scala 276:19]
  wire [29:0] csr_io_pmp_0_addr; // @[RocketCore.scala 276:19]
  wire [31:0] csr_io_pmp_0_mask; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_1_cfg_l; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_pmp_1_cfg_a; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_1_cfg_x; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_1_cfg_w; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_1_cfg_r; // @[RocketCore.scala 276:19]
  wire [29:0] csr_io_pmp_1_addr; // @[RocketCore.scala 276:19]
  wire [31:0] csr_io_pmp_1_mask; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_2_cfg_l; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_pmp_2_cfg_a; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_2_cfg_x; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_2_cfg_w; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_2_cfg_r; // @[RocketCore.scala 276:19]
  wire [29:0] csr_io_pmp_2_addr; // @[RocketCore.scala 276:19]
  wire [31:0] csr_io_pmp_2_mask; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_3_cfg_l; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_pmp_3_cfg_a; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_3_cfg_x; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_3_cfg_w; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_3_cfg_r; // @[RocketCore.scala 276:19]
  wire [29:0] csr_io_pmp_3_addr; // @[RocketCore.scala 276:19]
  wire [31:0] csr_io_pmp_3_mask; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_4_cfg_l; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_pmp_4_cfg_a; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_4_cfg_x; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_4_cfg_w; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_4_cfg_r; // @[RocketCore.scala 276:19]
  wire [29:0] csr_io_pmp_4_addr; // @[RocketCore.scala 276:19]
  wire [31:0] csr_io_pmp_4_mask; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_5_cfg_l; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_pmp_5_cfg_a; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_5_cfg_x; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_5_cfg_w; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_5_cfg_r; // @[RocketCore.scala 276:19]
  wire [29:0] csr_io_pmp_5_addr; // @[RocketCore.scala 276:19]
  wire [31:0] csr_io_pmp_5_mask; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_6_cfg_l; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_pmp_6_cfg_a; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_6_cfg_x; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_6_cfg_w; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_6_cfg_r; // @[RocketCore.scala 276:19]
  wire [29:0] csr_io_pmp_6_addr; // @[RocketCore.scala 276:19]
  wire [31:0] csr_io_pmp_6_mask; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_7_cfg_l; // @[RocketCore.scala 276:19]
  wire [1:0] csr_io_pmp_7_cfg_a; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_7_cfg_x; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_7_cfg_w; // @[RocketCore.scala 276:19]
  wire  csr_io_pmp_7_cfg_r; // @[RocketCore.scala 276:19]
  wire [29:0] csr_io_pmp_7_addr; // @[RocketCore.scala 276:19]
  wire [31:0] csr_io_pmp_7_mask; // @[RocketCore.scala 276:19]
  wire [31:0] csr_io_inst_0; // @[RocketCore.scala 276:19]
  wire  csr_io_trace_0_valid; // @[RocketCore.scala 276:19]
  wire [39:0] csr_io_trace_0_iaddr; // @[RocketCore.scala 276:19]
  wire [31:0] csr_io_trace_0_insn; // @[RocketCore.scala 276:19]
  wire  csr_io_trace_0_exception; // @[RocketCore.scala 276:19]
  wire [63:0] csr_io_customCSRs_0_value; // @[RocketCore.scala 276:19]
  wire [29:0] csr_io_covSum; // @[RocketCore.scala 276:19]
  wire  csr_metaAssert; // @[RocketCore.scala 276:19]
  wire  csr_metaReset; // @[RocketCore.scala 276:19]
  wire  bpu_io_status_debug; // @[RocketCore.scala 317:19]
  wire [1:0] bpu_io_status_prv; // @[RocketCore.scala 317:19]
  wire  bpu_io_bp_0_control_action; // @[RocketCore.scala 317:19]
  wire [1:0] bpu_io_bp_0_control_tmatch; // @[RocketCore.scala 317:19]
  wire  bpu_io_bp_0_control_m; // @[RocketCore.scala 317:19]
  wire  bpu_io_bp_0_control_s; // @[RocketCore.scala 317:19]
  wire  bpu_io_bp_0_control_u; // @[RocketCore.scala 317:19]
  wire  bpu_io_bp_0_control_x; // @[RocketCore.scala 317:19]
  wire  bpu_io_bp_0_control_w; // @[RocketCore.scala 317:19]
  wire  bpu_io_bp_0_control_r; // @[RocketCore.scala 317:19]
  wire [38:0] bpu_io_bp_0_address; // @[RocketCore.scala 317:19]
  wire [38:0] bpu_io_pc; // @[RocketCore.scala 317:19]
  wire [38:0] bpu_io_ea; // @[RocketCore.scala 317:19]
  wire  bpu_io_xcpt_if; // @[RocketCore.scala 317:19]
  wire  bpu_io_xcpt_ld; // @[RocketCore.scala 317:19]
  wire  bpu_io_xcpt_st; // @[RocketCore.scala 317:19]
  wire  bpu_io_debug_if; // @[RocketCore.scala 317:19]
  wire  bpu_io_debug_ld; // @[RocketCore.scala 317:19]
  wire  bpu_io_debug_st; // @[RocketCore.scala 317:19]
  wire [29:0] bpu_io_covSum; // @[RocketCore.scala 317:19]
  wire  bpu_metaAssert; // @[RocketCore.scala 317:19]
  wire  alu_io_dw; // @[RocketCore.scala 377:19]
  wire [3:0] alu_io_fn; // @[RocketCore.scala 377:19]
  wire [63:0] alu_io_in2; // @[RocketCore.scala 377:19]
  wire [63:0] alu_io_in1; // @[RocketCore.scala 377:19]
  wire [63:0] alu_io_out; // @[RocketCore.scala 377:19]
  wire [63:0] alu_io_adder_out; // @[RocketCore.scala 377:19]
  wire  alu_io_cmp_out; // @[RocketCore.scala 377:19]
  wire [29:0] alu_io_covSum; // @[RocketCore.scala 377:19]
  wire  alu_metaAssert; // @[RocketCore.scala 377:19]
  wire  div_clock; // @[RocketCore.scala 401:19]
  wire  div_reset; // @[RocketCore.scala 401:19]
  wire  div_io_req_ready; // @[RocketCore.scala 401:19]
  wire  div_io_req_valid; // @[RocketCore.scala 401:19]
  wire [3:0] div_io_req_bits_fn; // @[RocketCore.scala 401:19]
  wire  div_io_req_bits_dw; // @[RocketCore.scala 401:19]
  wire [63:0] div_io_req_bits_in1; // @[RocketCore.scala 401:19]
  wire [63:0] div_io_req_bits_in2; // @[RocketCore.scala 401:19]
  wire [4:0] div_io_req_bits_tag; // @[RocketCore.scala 401:19]
  wire  div_io_kill; // @[RocketCore.scala 401:19]
  wire  div_io_resp_ready; // @[RocketCore.scala 401:19]
  wire  div_io_resp_valid; // @[RocketCore.scala 401:19]
  wire [63:0] div_io_resp_bits_data; // @[RocketCore.scala 401:19]
  wire [4:0] div_io_resp_bits_tag; // @[RocketCore.scala 401:19]
  wire [29:0] div_io_covSum; // @[RocketCore.scala 401:19]
  wire  div_metaAssert; // @[RocketCore.scala 401:19]
  wire  div_metaReset; // @[RocketCore.scala 401:19]
  wire [29:0] PlusArgTimeout_io_covSum; // @[PlusArg.scala 89:11]
  wire  PlusArgTimeout_metaAssert; // @[PlusArg.scala 89:11]
  reg  id_reg_pause; // @[RocketCore.scala 110:25]
  reg [31:0] _RAND_3;
  reg  imem_might_request_reg; // @[RocketCore.scala 111:35]
  reg [31:0] _RAND_4;
  reg  ex_ctrl_fp; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_5;
  reg  ex_ctrl_branch; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_6;
  reg  ex_ctrl_jal; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_7;
  reg  ex_ctrl_jalr; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_8;
  reg  ex_ctrl_rxs2; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_9;
  reg  ex_ctrl_rxs1; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_10;
  reg [1:0] ex_ctrl_sel_alu2; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_11;
  reg [1:0] ex_ctrl_sel_alu1; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_12;
  reg [2:0] ex_ctrl_sel_imm; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_13;
  reg  ex_ctrl_alu_dw; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_14;
  reg [3:0] ex_ctrl_alu_fn; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_15;
  reg  ex_ctrl_mem; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_16;
  reg [4:0] ex_ctrl_mem_cmd; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_17;
  reg  ex_ctrl_rfs1; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_18;
  reg  ex_ctrl_rfs2; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_19;
  reg  ex_ctrl_wfd; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_20;
  reg  ex_ctrl_div; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_21;
  reg  ex_ctrl_wxd; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_22;
  reg [2:0] ex_ctrl_csr; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_23;
  reg  ex_ctrl_fence_i; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_24;
  reg  mem_ctrl_fp; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_25;
  reg  mem_ctrl_branch; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_26;
  reg  mem_ctrl_jal; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_27;
  reg  mem_ctrl_jalr; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_28;
  reg  mem_ctrl_rxs2; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_29;
  reg  mem_ctrl_rxs1; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_30;
  reg  mem_ctrl_mem; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_31;
  reg  mem_ctrl_rfs1; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_32;
  reg  mem_ctrl_rfs2; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_33;
  reg  mem_ctrl_wfd; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_34;
  reg  mem_ctrl_div; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_35;
  reg  mem_ctrl_wxd; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_36;
  reg [2:0] mem_ctrl_csr; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_37;
  reg  mem_ctrl_fence_i; // @[RocketCore.scala 185:21]
  reg [31:0] _RAND_38;
  reg  wb_ctrl_rxs2; // @[RocketCore.scala 186:20]
  reg [31:0] _RAND_39;
  reg  wb_ctrl_rxs1; // @[RocketCore.scala 186:20]
  reg [31:0] _RAND_40;
  reg  wb_ctrl_mem; // @[RocketCore.scala 186:20]
  reg [31:0] _RAND_41;
  reg  wb_ctrl_rfs1; // @[RocketCore.scala 186:20]
  reg [31:0] _RAND_42;
  reg  wb_ctrl_rfs2; // @[RocketCore.scala 186:20]
  reg [31:0] _RAND_43;
  reg  wb_ctrl_wfd; // @[RocketCore.scala 186:20]
  reg [31:0] _RAND_44;
  reg  wb_ctrl_div; // @[RocketCore.scala 186:20]
  reg [31:0] _RAND_45;
  reg  wb_ctrl_wxd; // @[RocketCore.scala 186:20]
  reg [31:0] _RAND_46;
  reg [2:0] wb_ctrl_csr; // @[RocketCore.scala 186:20]
  reg [31:0] _RAND_47;
  reg  wb_ctrl_fence_i; // @[RocketCore.scala 186:20]
  reg [31:0] _RAND_48;
  reg  ex_reg_xcpt_interrupt; // @[RocketCore.scala 188:35]
  reg [31:0] _RAND_49;
  reg  ex_reg_valid; // @[RocketCore.scala 189:35]
  reg [31:0] _RAND_50;
  reg  ex_reg_rvc; // @[RocketCore.scala 190:35]
  reg [31:0] _RAND_51;
  reg [4:0] ex_reg_btb_resp_entry; // @[RocketCore.scala 191:35]
  reg [31:0] _RAND_52;
  reg [7:0] ex_reg_btb_resp_bht_history; // @[RocketCore.scala 191:35]
  reg [31:0] _RAND_53;
  reg  ex_reg_xcpt; // @[RocketCore.scala 192:35]
  reg [31:0] _RAND_54;
  reg  ex_reg_flush_pipe; // @[RocketCore.scala 193:35]
  reg [31:0] _RAND_55;
  reg  ex_reg_load_use; // @[RocketCore.scala 194:35]
  reg [31:0] _RAND_56;
  reg [63:0] ex_reg_cause; // @[RocketCore.scala 195:35]
  reg [63:0] _RAND_57;
  reg  ex_reg_replay; // @[RocketCore.scala 196:26]
  reg [31:0] _RAND_58;
  reg [39:0] ex_reg_pc; // @[RocketCore.scala 197:22]
  reg [63:0] _RAND_59;
  reg [1:0] ex_reg_mem_size; // @[RocketCore.scala 198:28]
  reg [31:0] _RAND_60;
  reg [31:0] ex_reg_inst; // @[RocketCore.scala 199:24]
  reg [31:0] _RAND_61;
  reg [31:0] ex_reg_raw_inst; // @[RocketCore.scala 200:28]
  reg [31:0] _RAND_62;
  reg  mem_reg_xcpt_interrupt; // @[RocketCore.scala 205:36]
  reg [31:0] _RAND_63;
  reg  mem_reg_valid; // @[RocketCore.scala 206:36]
  reg [31:0] _RAND_64;
  reg  mem_reg_rvc; // @[RocketCore.scala 207:36]
  reg [31:0] _RAND_65;
  reg [4:0] mem_reg_btb_resp_entry; // @[RocketCore.scala 208:36]
  reg [31:0] _RAND_66;
  reg [7:0] mem_reg_btb_resp_bht_history; // @[RocketCore.scala 208:36]
  reg [31:0] _RAND_67;
  reg  mem_reg_xcpt; // @[RocketCore.scala 209:36]
  reg [31:0] _RAND_68;
  reg  mem_reg_replay; // @[RocketCore.scala 210:36]
  reg [31:0] _RAND_69;
  reg  mem_reg_flush_pipe; // @[RocketCore.scala 211:36]
  reg [31:0] _RAND_70;
  reg [63:0] mem_reg_cause; // @[RocketCore.scala 212:36]
  reg [63:0] _RAND_71;
  reg  mem_reg_slow_bypass; // @[RocketCore.scala 213:36]
  reg [31:0] _RAND_72;
  reg  mem_reg_load; // @[RocketCore.scala 214:36]
  reg [31:0] _RAND_73;
  reg  mem_reg_store; // @[RocketCore.scala 215:36]
  reg [31:0] _RAND_74;
  reg  mem_reg_sfence; // @[RocketCore.scala 216:27]
  reg [31:0] _RAND_75;
  reg [39:0] mem_reg_pc; // @[RocketCore.scala 217:23]
  reg [63:0] _RAND_76;
  reg [31:0] mem_reg_inst; // @[RocketCore.scala 218:25]
  reg [31:0] _RAND_77;
  reg [1:0] mem_reg_mem_size; // @[RocketCore.scala 219:29]
  reg [31:0] _RAND_78;
  reg [31:0] mem_reg_raw_inst; // @[RocketCore.scala 220:29]
  reg [31:0] _RAND_79;
  reg [63:0] mem_reg_wdata; // @[RocketCore.scala 223:26]
  reg [63:0] _RAND_80;
  reg [63:0] mem_reg_rs2; // @[RocketCore.scala 224:24]
  reg [63:0] _RAND_81;
  reg  mem_br_taken; // @[RocketCore.scala 225:25]
  reg [31:0] _RAND_82;
  reg  wb_reg_valid; // @[RocketCore.scala 229:35]
  reg [31:0] _RAND_83;
  reg  wb_reg_xcpt; // @[RocketCore.scala 230:35]
  reg [31:0] _RAND_84;
  reg  wb_reg_replay; // @[RocketCore.scala 231:35]
  reg [31:0] _RAND_85;
  reg  wb_reg_flush_pipe; // @[RocketCore.scala 232:35]
  reg [31:0] _RAND_86;
  reg [63:0] wb_reg_cause; // @[RocketCore.scala 233:35]
  reg [63:0] _RAND_87;
  reg  wb_reg_sfence; // @[RocketCore.scala 234:26]
  reg [31:0] _RAND_88;
  reg [39:0] wb_reg_pc; // @[RocketCore.scala 235:22]
  reg [63:0] _RAND_89;
  reg [1:0] wb_reg_mem_size; // @[RocketCore.scala 236:28]
  reg [31:0] _RAND_90;
  reg [31:0] wb_reg_inst; // @[RocketCore.scala 237:24]
  reg [31:0] _RAND_91;
  reg [31:0] wb_reg_raw_inst; // @[RocketCore.scala 238:28]
  reg [31:0] _RAND_92;
  reg [63:0] wb_reg_wdata; // @[RocketCore.scala 239:25]
  reg [63:0] _RAND_93;
  wire  replay_wb_common; // @[RocketCore.scala 629:42]
  wire  _T_1465; // @[RocketCore.scala 607:19]
  wire  _T_1466; // @[RocketCore.scala 607:34]
  wire  _T_1477; // @[RocketCore.scala 974:26]
  wire  _T_1468; // @[RocketCore.scala 608:34]
  wire  _T_1478; // @[RocketCore.scala 974:26]
  wire  _T_1470; // @[RocketCore.scala 609:34]
  wire  _T_1479; // @[RocketCore.scala 974:26]
  wire  _T_1472; // @[RocketCore.scala 610:34]
  wire  _T_1480; // @[RocketCore.scala 974:26]
  wire  _T_1474; // @[RocketCore.scala 611:34]
  wire  _T_1481; // @[RocketCore.scala 974:26]
  wire  _T_1476; // @[RocketCore.scala 612:34]
  wire  wb_xcpt; // @[RocketCore.scala 974:26]
  wire  _T_1503; // @[RocketCore.scala 632:27]
  wire  _T_1504; // @[RocketCore.scala 632:38]
  wire  take_pc_wb; // @[RocketCore.scala 632:53]
  wire  _T_1149; // @[RocketCore.scala 482:34]
  wire  ex_pc_valid; // @[RocketCore.scala 482:51]
  wire  _T_1305; // @[RocketCore.scala 505:36]
  wire [24:0] a; // @[RocketCore.scala 988:23]
  wire  _T_1307; // @[RocketCore.scala 989:21]
  wire  _T_1308; // @[RocketCore.scala 989:34]
  wire  _T_1309; // @[RocketCore.scala 989:29]
  wire  msb; // @[RocketCore.scala 989:18]
  wire [39:0] _T_1315; // @[RocketCore.scala 505:106]
  wire  _T_1175; // @[RocketCore.scala 502:25]
  wire  _T_1178; // @[RocketCore.scala 1036:53]
  wire  _T_1233; // @[Cat.scala 29:58]
  wire [10:0] _T_1232; // @[Cat.scala 29:58]
  wire [7:0] _T_1230; // @[Cat.scala 29:58]
  wire  _T_1229; // @[Cat.scala 29:58]
  wire [31:0] _T_1237; // @[RocketCore.scala 1050:53]
  wire [7:0] _T_1292; // @[Cat.scala 29:58]
  wire  _T_1291; // @[Cat.scala 29:58]
  wire [31:0] _T_1299; // @[RocketCore.scala 1050:53]
  wire [3:0] _T_1300; // @[RocketCore.scala 504:8]
  wire [31:0] _T_1301; // @[RocketCore.scala 503:8]
  wire [31:0] _T_1302; // @[RocketCore.scala 502:8]
  wire [39:0] _GEN_248; // @[RocketCore.scala 501:41]
  wire [39:0] mem_br_target; // @[RocketCore.scala 501:41]
  wire [39:0] _T_1316; // @[RocketCore.scala 505:21]
  wire [39:0] mem_npc; // @[RocketCore.scala 505:141]
  wire  _T_1319; // @[RocketCore.scala 507:30]
  wire  _T_1320; // @[RocketCore.scala 508:31]
  wire  _T_1321; // @[RocketCore.scala 508:62]
  wire  _T_1322; // @[RocketCore.scala 508:8]
  wire  mem_wrong_npc; // @[RocketCore.scala 507:8]
  wire  _T_1338; // @[RocketCore.scala 515:54]
  wire  take_pc_mem; // @[RocketCore.scala 515:32]
  wire  take_pc_mem_wb; // @[RocketCore.scala 244:35]
  wire [31:0] _T_3; // @[Decode.scala 14:65]
  wire  _T_4; // @[Decode.scala 14:121]
  wire  _T_6; // @[Decode.scala 14:121]
  wire  _T_8; // @[Decode.scala 14:121]
  wire  _T_10; // @[Decode.scala 14:121]
  wire  _T_12; // @[Decode.scala 14:121]
  wire  _T_14; // @[Decode.scala 14:121]
  wire  _T_16; // @[Decode.scala 14:121]
  wire  _T_18; // @[Decode.scala 14:121]
  wire  _T_20; // @[Decode.scala 14:121]
  wire  _T_22; // @[Decode.scala 14:121]
  wire  _T_24; // @[Decode.scala 14:121]
  wire  _T_26; // @[Decode.scala 14:121]
  wire  _T_28; // @[Decode.scala 14:121]
  wire [31:0] _T_29; // @[Decode.scala 14:65]
  wire  _T_30; // @[Decode.scala 14:121]
  wire  _T_32; // @[Decode.scala 14:121]
  wire  _T_34; // @[Decode.scala 14:121]
  wire  _T_36; // @[Decode.scala 14:121]
  wire  _T_38; // @[Decode.scala 14:121]
  wire  _T_40; // @[Decode.scala 14:121]
  wire  _T_42; // @[Decode.scala 14:121]
  wire  _T_44; // @[Decode.scala 14:121]
  wire  _T_46; // @[Decode.scala 14:121]
  wire [31:0] _T_47; // @[Decode.scala 14:65]
  wire  _T_48; // @[Decode.scala 14:121]
  wire  _T_50; // @[Decode.scala 14:121]
  wire  _T_52; // @[Decode.scala 14:121]
  wire  _T_54; // @[Decode.scala 14:121]
  wire  _T_56; // @[Decode.scala 14:121]
  wire  _T_58; // @[Decode.scala 14:121]
  wire  _T_60; // @[Decode.scala 14:121]
  wire  _T_62; // @[Decode.scala 14:121]
  wire  _T_64; // @[Decode.scala 14:121]
  wire  _T_66; // @[Decode.scala 14:121]
  wire  _T_68; // @[Decode.scala 14:121]
  wire  _T_70; // @[Decode.scala 14:121]
  wire  _T_72; // @[Decode.scala 14:121]
  wire  _T_74; // @[Decode.scala 14:121]
  wire  _T_76; // @[Decode.scala 14:121]
  wire  _T_78; // @[Decode.scala 14:121]
  wire  _T_80; // @[Decode.scala 14:121]
  wire  _T_82; // @[Decode.scala 14:121]
  wire [31:0] _T_83; // @[Decode.scala 14:65]
  wire  _T_84; // @[Decode.scala 14:121]
  wire  _T_86; // @[Decode.scala 14:121]
  wire  _T_88; // @[Decode.scala 14:121]
  wire [31:0] _T_89; // @[Decode.scala 14:65]
  wire  _T_90; // @[Decode.scala 14:121]
  wire  _T_92; // @[Decode.scala 14:121]
  wire  _T_94; // @[Decode.scala 14:121]
  wire  _T_96; // @[Decode.scala 14:121]
  wire [31:0] _T_97; // @[Decode.scala 14:65]
  wire  _T_98; // @[Decode.scala 14:121]
  wire  _T_100; // @[Decode.scala 14:121]
  wire [31:0] _T_101; // @[Decode.scala 14:65]
  wire  _T_102; // @[Decode.scala 14:121]
  wire  _T_104; // @[Decode.scala 14:121]
  wire  _T_106; // @[Decode.scala 14:121]
  wire  _T_108; // @[Decode.scala 14:121]
  wire  _T_110; // @[Decode.scala 14:121]
  wire  _T_112; // @[Decode.scala 14:121]
  wire  _T_114; // @[Decode.scala 14:121]
  wire  _T_116; // @[Decode.scala 14:121]
  wire [31:0] _T_117; // @[Decode.scala 14:65]
  wire  _T_118; // @[Decode.scala 14:121]
  wire  _T_120; // @[Decode.scala 14:121]
  wire  _T_122; // @[Decode.scala 14:121]
  wire  _T_124; // @[Decode.scala 14:121]
  wire  _T_126; // @[Decode.scala 14:121]
  wire  _T_128; // @[Decode.scala 14:121]
  wire  _T_130; // @[Decode.scala 14:121]
  wire  _T_132; // @[Decode.scala 14:121]
  wire  _T_134; // @[Decode.scala 14:121]
  wire  _T_136; // @[Decode.scala 14:121]
  wire  _T_138; // @[Decode.scala 14:121]
  wire  _T_140; // @[Decode.scala 14:121]
  wire  _T_142; // @[Decode.scala 14:121]
  wire  _T_144; // @[Decode.scala 14:121]
  wire  _T_146; // @[Decode.scala 14:121]
  wire  _T_148; // @[Decode.scala 14:121]
  wire  _T_150; // @[Decode.scala 14:121]
  wire  _T_152; // @[Decode.scala 14:121]
  wire  _T_154; // @[Decode.scala 14:121]
  wire  _T_156; // @[Decode.scala 14:121]
  wire  _T_158; // @[Decode.scala 14:121]
  wire  _T_160; // @[Decode.scala 14:121]
  wire  _T_162; // @[Decode.scala 14:121]
  wire  _T_164; // @[Decode.scala 14:121]
  wire  _T_166; // @[Decode.scala 14:121]
  wire  _T_168; // @[Decode.scala 14:121]
  wire  _T_170; // @[Decode.scala 14:121]
  wire  _T_172; // @[Decode.scala 14:121]
  wire  _T_174; // @[Decode.scala 14:121]
  wire  _T_176; // @[Decode.scala 14:121]
  wire  _T_178; // @[Decode.scala 14:121]
  wire  _T_180; // @[Decode.scala 14:121]
  wire  _T_182; // @[Decode.scala 14:121]
  wire  _T_184; // @[Decode.scala 14:121]
  wire  _T_186; // @[Decode.scala 14:121]
  wire  _T_188; // @[Decode.scala 14:121]
  wire  _T_190; // @[Decode.scala 14:121]
  wire  _T_192; // @[Decode.scala 14:121]
  wire  _T_194; // @[Decode.scala 14:121]
  wire  _T_196; // @[Decode.scala 14:121]
  wire  _T_198; // @[Decode.scala 14:121]
  wire  _T_200; // @[Decode.scala 14:121]
  wire  _T_202; // @[Decode.scala 14:121]
  wire [31:0] _T_203; // @[Decode.scala 14:65]
  wire  _T_204; // @[Decode.scala 14:121]
  wire  _T_206; // @[Decode.scala 14:121]
  wire  _T_208; // @[Decode.scala 14:121]
  wire  _T_210; // @[Decode.scala 14:121]
  wire  _T_212; // @[Decode.scala 14:121]
  wire  _T_214; // @[Decode.scala 14:121]
  wire  _T_216; // @[Decode.scala 14:121]
  wire  _T_218; // @[Decode.scala 14:121]
  wire  _T_220; // @[Decode.scala 14:121]
  wire  _T_222; // @[Decode.scala 14:121]
  wire  _T_224; // @[Decode.scala 14:121]
  wire  _T_226; // @[Decode.scala 14:121]
  wire [31:0] _T_227; // @[Decode.scala 14:65]
  wire  _T_228; // @[Decode.scala 14:121]
  wire  _T_229; // @[Decode.scala 14:121]
  wire  _T_230; // @[Decode.scala 14:121]
  wire  _T_232; // @[Decode.scala 14:121]
  wire  _T_234; // @[Decode.scala 14:121]
  wire  _T_236; // @[Decode.scala 14:121]
  wire  _T_238; // @[Decode.scala 14:121]
  wire  _T_240; // @[Decode.scala 14:121]
  wire  _T_242; // @[Decode.scala 14:121]
  wire  _T_244; // @[Decode.scala 14:121]
  wire [31:0] _T_245; // @[Decode.scala 14:65]
  wire  _T_246; // @[Decode.scala 14:121]
  wire  _T_248; // @[Decode.scala 14:121]
  wire  _T_250; // @[Decode.scala 14:121]
  wire  _T_252; // @[Decode.scala 14:121]
  wire  _T_254; // @[Decode.scala 14:121]
  wire  _T_256; // @[Decode.scala 14:121]
  wire  _T_258; // @[Decode.scala 14:121]
  wire  _T_260; // @[Decode.scala 14:121]
  wire  _T_262; // @[Decode.scala 14:121]
  wire  _T_264; // @[Decode.scala 14:121]
  wire  _T_266; // @[Decode.scala 14:121]
  wire  _T_268; // @[Decode.scala 14:121]
  wire  _T_270; // @[Decode.scala 14:121]
  wire  _T_272; // @[Decode.scala 14:121]
  wire  _T_274; // @[Decode.scala 14:121]
  wire  _T_276; // @[Decode.scala 14:121]
  wire  _T_278; // @[Decode.scala 14:121]
  wire  _T_280; // @[Decode.scala 14:121]
  wire  _T_282; // @[Decode.scala 14:121]
  wire  _T_284; // @[Decode.scala 14:121]
  wire  _T_286; // @[Decode.scala 14:121]
  wire  _T_288; // @[Decode.scala 14:121]
  wire  _T_290; // @[Decode.scala 14:121]
  wire  _T_292; // @[Decode.scala 14:121]
  wire  _T_294; // @[Decode.scala 14:121]
  wire  _T_296; // @[Decode.scala 14:121]
  wire  _T_298; // @[Decode.scala 14:121]
  wire  _T_300; // @[Decode.scala 14:121]
  wire  _T_302; // @[Decode.scala 14:121]
  wire  _T_303; // @[Decode.scala 14:121]
  wire  _T_304; // @[Decode.scala 14:121]
  wire  _T_305; // @[Decode.scala 14:121]
  wire  _T_306; // @[Decode.scala 14:121]
  wire  _T_307; // @[Decode.scala 14:121]
  wire  _T_309; // @[Decode.scala 14:121]
  wire  _T_311; // @[Decode.scala 14:121]
  wire  _T_313; // @[Decode.scala 14:121]
  wire  _T_315; // @[Decode.scala 14:121]
  wire  _T_317; // @[Decode.scala 14:121]
  wire  _T_319; // @[Decode.scala 14:121]
  wire  _T_321; // @[Decode.scala 15:30]
  wire  _T_322; // @[Decode.scala 15:30]
  wire  _T_323; // @[Decode.scala 15:30]
  wire  _T_324; // @[Decode.scala 15:30]
  wire  _T_325; // @[Decode.scala 15:30]
  wire  _T_326; // @[Decode.scala 15:30]
  wire  _T_327; // @[Decode.scala 15:30]
  wire  _T_328; // @[Decode.scala 15:30]
  wire  _T_329; // @[Decode.scala 15:30]
  wire  _T_330; // @[Decode.scala 15:30]
  wire  _T_331; // @[Decode.scala 15:30]
  wire  _T_332; // @[Decode.scala 15:30]
  wire  _T_333; // @[Decode.scala 15:30]
  wire  _T_334; // @[Decode.scala 15:30]
  wire  _T_335; // @[Decode.scala 15:30]
  wire  _T_336; // @[Decode.scala 15:30]
  wire  _T_337; // @[Decode.scala 15:30]
  wire  _T_338; // @[Decode.scala 15:30]
  wire  _T_339; // @[Decode.scala 15:30]
  wire  _T_340; // @[Decode.scala 15:30]
  wire  _T_341; // @[Decode.scala 15:30]
  wire  _T_342; // @[Decode.scala 15:30]
  wire  _T_343; // @[Decode.scala 15:30]
  wire  _T_344; // @[Decode.scala 15:30]
  wire  _T_345; // @[Decode.scala 15:30]
  wire  _T_346; // @[Decode.scala 15:30]
  wire  _T_347; // @[Decode.scala 15:30]
  wire  _T_348; // @[Decode.scala 15:30]
  wire  _T_349; // @[Decode.scala 15:30]
  wire  _T_350; // @[Decode.scala 15:30]
  wire  _T_351; // @[Decode.scala 15:30]
  wire  _T_352; // @[Decode.scala 15:30]
  wire  _T_353; // @[Decode.scala 15:30]
  wire  _T_354; // @[Decode.scala 15:30]
  wire  _T_355; // @[Decode.scala 15:30]
  wire  _T_356; // @[Decode.scala 15:30]
  wire  _T_357; // @[Decode.scala 15:30]
  wire  _T_358; // @[Decode.scala 15:30]
  wire  _T_359; // @[Decode.scala 15:30]
  wire  _T_360; // @[Decode.scala 15:30]
  wire  _T_361; // @[Decode.scala 15:30]
  wire  _T_362; // @[Decode.scala 15:30]
  wire  _T_363; // @[Decode.scala 15:30]
  wire  _T_364; // @[Decode.scala 15:30]
  wire  _T_365; // @[Decode.scala 15:30]
  wire  _T_366; // @[Decode.scala 15:30]
  wire  _T_367; // @[Decode.scala 15:30]
  wire  _T_368; // @[Decode.scala 15:30]
  wire  _T_369; // @[Decode.scala 15:30]
  wire  _T_370; // @[Decode.scala 15:30]
  wire  _T_371; // @[Decode.scala 15:30]
  wire  _T_372; // @[Decode.scala 15:30]
  wire  _T_373; // @[Decode.scala 15:30]
  wire  _T_374; // @[Decode.scala 15:30]
  wire  _T_375; // @[Decode.scala 15:30]
  wire  _T_376; // @[Decode.scala 15:30]
  wire  _T_377; // @[Decode.scala 15:30]
  wire  _T_378; // @[Decode.scala 15:30]
  wire  _T_379; // @[Decode.scala 15:30]
  wire  _T_380; // @[Decode.scala 15:30]
  wire  _T_381; // @[Decode.scala 15:30]
  wire  _T_382; // @[Decode.scala 15:30]
  wire  _T_383; // @[Decode.scala 15:30]
  wire  _T_384; // @[Decode.scala 15:30]
  wire  _T_385; // @[Decode.scala 15:30]
  wire  _T_386; // @[Decode.scala 15:30]
  wire  _T_387; // @[Decode.scala 15:30]
  wire  _T_388; // @[Decode.scala 15:30]
  wire  _T_389; // @[Decode.scala 15:30]
  wire  _T_390; // @[Decode.scala 15:30]
  wire  _T_391; // @[Decode.scala 15:30]
  wire  _T_392; // @[Decode.scala 15:30]
  wire  _T_393; // @[Decode.scala 15:30]
  wire  _T_394; // @[Decode.scala 15:30]
  wire  _T_395; // @[Decode.scala 15:30]
  wire  _T_396; // @[Decode.scala 15:30]
  wire  _T_397; // @[Decode.scala 15:30]
  wire  _T_398; // @[Decode.scala 15:30]
  wire  _T_399; // @[Decode.scala 15:30]
  wire  _T_400; // @[Decode.scala 15:30]
  wire  _T_401; // @[Decode.scala 15:30]
  wire  _T_402; // @[Decode.scala 15:30]
  wire  _T_403; // @[Decode.scala 15:30]
  wire  _T_404; // @[Decode.scala 15:30]
  wire  _T_405; // @[Decode.scala 15:30]
  wire  _T_406; // @[Decode.scala 15:30]
  wire  _T_407; // @[Decode.scala 15:30]
  wire  _T_408; // @[Decode.scala 15:30]
  wire  _T_409; // @[Decode.scala 15:30]
  wire  _T_410; // @[Decode.scala 15:30]
  wire  _T_411; // @[Decode.scala 15:30]
  wire  _T_412; // @[Decode.scala 15:30]
  wire  _T_413; // @[Decode.scala 15:30]
  wire  _T_414; // @[Decode.scala 15:30]
  wire  _T_415; // @[Decode.scala 15:30]
  wire  _T_416; // @[Decode.scala 15:30]
  wire  _T_417; // @[Decode.scala 15:30]
  wire  _T_418; // @[Decode.scala 15:30]
  wire  _T_419; // @[Decode.scala 15:30]
  wire  _T_420; // @[Decode.scala 15:30]
  wire  _T_421; // @[Decode.scala 15:30]
  wire  _T_422; // @[Decode.scala 15:30]
  wire  _T_423; // @[Decode.scala 15:30]
  wire  _T_424; // @[Decode.scala 15:30]
  wire  _T_425; // @[Decode.scala 15:30]
  wire  _T_426; // @[Decode.scala 15:30]
  wire  _T_427; // @[Decode.scala 15:30]
  wire  _T_428; // @[Decode.scala 15:30]
  wire  _T_429; // @[Decode.scala 15:30]
  wire  _T_430; // @[Decode.scala 15:30]
  wire  _T_431; // @[Decode.scala 15:30]
  wire  _T_432; // @[Decode.scala 15:30]
  wire  _T_433; // @[Decode.scala 15:30]
  wire  _T_434; // @[Decode.scala 15:30]
  wire  _T_435; // @[Decode.scala 15:30]
  wire  _T_436; // @[Decode.scala 15:30]
  wire  _T_437; // @[Decode.scala 15:30]
  wire  _T_438; // @[Decode.scala 15:30]
  wire  _T_439; // @[Decode.scala 15:30]
  wire  _T_440; // @[Decode.scala 15:30]
  wire  _T_441; // @[Decode.scala 15:30]
  wire  _T_442; // @[Decode.scala 15:30]
  wire  _T_443; // @[Decode.scala 15:30]
  wire  _T_444; // @[Decode.scala 15:30]
  wire  _T_445; // @[Decode.scala 15:30]
  wire  _T_446; // @[Decode.scala 15:30]
  wire  _T_447; // @[Decode.scala 15:30]
  wire  _T_448; // @[Decode.scala 15:30]
  wire  _T_449; // @[Decode.scala 15:30]
  wire  _T_450; // @[Decode.scala 15:30]
  wire  _T_451; // @[Decode.scala 15:30]
  wire  _T_452; // @[Decode.scala 15:30]
  wire  _T_453; // @[Decode.scala 15:30]
  wire  _T_454; // @[Decode.scala 15:30]
  wire  _T_455; // @[Decode.scala 15:30]
  wire  _T_456; // @[Decode.scala 15:30]
  wire  _T_457; // @[Decode.scala 15:30]
  wire  _T_458; // @[Decode.scala 15:30]
  wire  _T_459; // @[Decode.scala 15:30]
  wire  _T_460; // @[Decode.scala 15:30]
  wire  _T_461; // @[Decode.scala 15:30]
  wire  _T_462; // @[Decode.scala 15:30]
  wire  _T_463; // @[Decode.scala 15:30]
  wire  _T_464; // @[Decode.scala 15:30]
  wire  _T_465; // @[Decode.scala 15:30]
  wire  _T_466; // @[Decode.scala 15:30]
  wire  _T_467; // @[Decode.scala 15:30]
  wire  _T_468; // @[Decode.scala 15:30]
  wire  _T_469; // @[Decode.scala 15:30]
  wire  _T_470; // @[Decode.scala 15:30]
  wire  _T_471; // @[Decode.scala 15:30]
  wire  _T_472; // @[Decode.scala 15:30]
  wire  _T_473; // @[Decode.scala 15:30]
  wire  _T_474; // @[Decode.scala 15:30]
  wire  _T_475; // @[Decode.scala 15:30]
  wire  _T_476; // @[Decode.scala 15:30]
  wire  _T_477; // @[Decode.scala 15:30]
  wire  _T_478; // @[Decode.scala 15:30]
  wire  _T_479; // @[Decode.scala 15:30]
  wire  _T_480; // @[Decode.scala 15:30]
  wire  id_ctrl_legal; // @[Decode.scala 15:30]
  wire [31:0] _T_482; // @[Decode.scala 14:65]
  wire  _T_483; // @[Decode.scala 14:121]
  wire [31:0] _T_484; // @[Decode.scala 14:65]
  wire  _T_485; // @[Decode.scala 14:121]
  wire  id_ctrl_fp; // @[Decode.scala 15:30]
  wire [31:0] _T_488; // @[Decode.scala 14:65]
  wire  id_ctrl_branch; // @[Decode.scala 14:121]
  wire [31:0] _T_491; // @[Decode.scala 14:65]
  wire  id_ctrl_jal; // @[Decode.scala 14:121]
  wire [31:0] _T_494; // @[Decode.scala 14:65]
  wire  id_ctrl_jalr; // @[Decode.scala 14:121]
  wire [31:0] _T_497; // @[Decode.scala 14:65]
  wire  _T_498; // @[Decode.scala 14:121]
  wire [31:0] _T_499; // @[Decode.scala 14:65]
  wire  _T_500; // @[Decode.scala 14:121]
  wire [31:0] _T_501; // @[Decode.scala 14:65]
  wire  _T_502; // @[Decode.scala 14:121]
  wire [31:0] _T_503; // @[Decode.scala 14:65]
  wire  _T_504; // @[Decode.scala 14:121]
  wire  _T_506; // @[Decode.scala 15:30]
  wire  _T_507; // @[Decode.scala 15:30]
  wire  id_ctrl_rxs2; // @[Decode.scala 15:30]
  wire [31:0] _T_509; // @[Decode.scala 14:65]
  wire  _T_510; // @[Decode.scala 14:121]
  wire [31:0] _T_511; // @[Decode.scala 14:65]
  wire  _T_512; // @[Decode.scala 14:121]
  wire [31:0] _T_513; // @[Decode.scala 14:65]
  wire  _T_514; // @[Decode.scala 14:121]
  wire [31:0] _T_515; // @[Decode.scala 14:65]
  wire  _T_516; // @[Decode.scala 14:121]
  wire [31:0] _T_517; // @[Decode.scala 14:65]
  wire  _T_518; // @[Decode.scala 14:121]
  wire  _T_520; // @[Decode.scala 15:30]
  wire  _T_521; // @[Decode.scala 15:30]
  wire  _T_522; // @[Decode.scala 15:30]
  wire  id_ctrl_rxs1; // @[Decode.scala 15:30]
  wire [31:0] _T_524; // @[Decode.scala 14:65]
  wire  _T_525; // @[Decode.scala 14:121]
  wire [31:0] _T_526; // @[Decode.scala 14:65]
  wire  _T_527; // @[Decode.scala 14:121]
  wire [31:0] _T_528; // @[Decode.scala 14:65]
  wire  _T_529; // @[Decode.scala 14:121]
  wire [31:0] _T_530; // @[Decode.scala 14:65]
  wire  _T_531; // @[Decode.scala 14:121]
  wire [31:0] _T_532; // @[Decode.scala 14:65]
  wire  _T_533; // @[Decode.scala 14:121]
  wire  _T_535; // @[Decode.scala 15:30]
  wire  _T_536; // @[Decode.scala 15:30]
  wire  _T_537; // @[Decode.scala 15:30]
  wire  _T_538; // @[Decode.scala 15:30]
  wire  _T_540; // @[Decode.scala 14:121]
  wire [31:0] _T_541; // @[Decode.scala 14:65]
  wire  _T_542; // @[Decode.scala 14:121]
  wire [31:0] _T_543; // @[Decode.scala 14:65]
  wire  _T_544; // @[Decode.scala 14:121]
  wire  _T_546; // @[Decode.scala 15:30]
  wire  _T_547; // @[Decode.scala 15:30]
  wire  _T_548; // @[Decode.scala 15:30]
  wire [1:0] id_ctrl_sel_alu2; // @[Cat.scala 29:58]
  wire [31:0] _T_550; // @[Decode.scala 14:65]
  wire  _T_551; // @[Decode.scala 14:121]
  wire [31:0] _T_552; // @[Decode.scala 14:65]
  wire  _T_553; // @[Decode.scala 14:121]
  wire [31:0] _T_554; // @[Decode.scala 14:65]
  wire  _T_555; // @[Decode.scala 14:121]
  wire  _T_557; // @[Decode.scala 15:30]
  wire  _T_558; // @[Decode.scala 15:30]
  wire  _T_559; // @[Decode.scala 15:30]
  wire  _T_560; // @[Decode.scala 15:30]
  wire  _T_562; // @[Decode.scala 14:121]
  wire  _T_564; // @[Decode.scala 15:30]
  wire [1:0] id_ctrl_sel_alu1; // @[Cat.scala 29:58]
  wire  _T_567; // @[Decode.scala 14:121]
  wire  _T_569; // @[Decode.scala 14:121]
  wire  _T_571; // @[Decode.scala 15:30]
  wire [31:0] _T_572; // @[Decode.scala 14:65]
  wire  _T_573; // @[Decode.scala 14:121]
  wire  _T_575; // @[Decode.scala 15:30]
  wire [31:0] _T_576; // @[Decode.scala 14:65]
  wire  _T_577; // @[Decode.scala 14:121]
  wire [31:0] _T_578; // @[Decode.scala 14:65]
  wire  _T_579; // @[Decode.scala 14:121]
  wire  _T_581; // @[Decode.scala 14:121]
  wire  _T_583; // @[Decode.scala 15:30]
  wire  _T_584; // @[Decode.scala 15:30]
  wire [2:0] id_ctrl_sel_imm; // @[Cat.scala 29:58]
  wire [31:0] _T_587; // @[Decode.scala 14:65]
  wire  _T_588; // @[Decode.scala 14:121]
  wire [31:0] _T_589; // @[Decode.scala 14:65]
  wire  _T_590; // @[Decode.scala 14:121]
  wire  id_ctrl_alu_dw; // @[Decode.scala 15:30]
  wire [31:0] _T_593; // @[Decode.scala 14:65]
  wire  _T_594; // @[Decode.scala 14:121]
  wire [31:0] _T_595; // @[Decode.scala 14:65]
  wire  _T_596; // @[Decode.scala 14:121]
  wire [31:0] _T_597; // @[Decode.scala 14:65]
  wire  _T_598; // @[Decode.scala 14:121]
  wire [31:0] _T_599; // @[Decode.scala 14:65]
  wire  _T_600; // @[Decode.scala 14:121]
  wire  _T_602; // @[Decode.scala 15:30]
  wire  _T_603; // @[Decode.scala 15:30]
  wire  _T_604; // @[Decode.scala 15:30]
  wire [31:0] _T_605; // @[Decode.scala 14:65]
  wire  _T_606; // @[Decode.scala 14:121]
  wire [31:0] _T_607; // @[Decode.scala 14:65]
  wire  _T_608; // @[Decode.scala 14:121]
  wire  _T_610; // @[Decode.scala 14:121]
  wire [31:0] _T_611; // @[Decode.scala 14:65]
  wire  _T_612; // @[Decode.scala 14:121]
  wire [31:0] _T_613; // @[Decode.scala 14:65]
  wire  _T_614; // @[Decode.scala 14:121]
  wire [31:0] _T_615; // @[Decode.scala 14:65]
  wire  _T_616; // @[Decode.scala 14:121]
  wire [31:0] _T_617; // @[Decode.scala 14:65]
  wire  _T_618; // @[Decode.scala 14:121]
  wire  _T_620; // @[Decode.scala 15:30]
  wire  _T_621; // @[Decode.scala 15:30]
  wire  _T_622; // @[Decode.scala 15:30]
  wire  _T_623; // @[Decode.scala 15:30]
  wire  _T_624; // @[Decode.scala 15:30]
  wire  _T_625; // @[Decode.scala 15:30]
  wire [31:0] _T_626; // @[Decode.scala 14:65]
  wire  _T_627; // @[Decode.scala 14:121]
  wire [31:0] _T_628; // @[Decode.scala 14:65]
  wire  _T_629; // @[Decode.scala 14:121]
  wire [31:0] _T_630; // @[Decode.scala 14:65]
  wire  _T_631; // @[Decode.scala 14:121]
  wire [31:0] _T_632; // @[Decode.scala 14:65]
  wire  _T_633; // @[Decode.scala 14:121]
  wire [31:0] _T_634; // @[Decode.scala 14:65]
  wire  _T_635; // @[Decode.scala 14:121]
  wire  _T_637; // @[Decode.scala 15:30]
  wire  _T_638; // @[Decode.scala 15:30]
  wire  _T_639; // @[Decode.scala 15:30]
  wire  _T_640; // @[Decode.scala 15:30]
  wire [31:0] _T_641; // @[Decode.scala 14:65]
  wire  _T_642; // @[Decode.scala 14:121]
  wire [31:0] _T_643; // @[Decode.scala 14:65]
  wire  _T_644; // @[Decode.scala 14:121]
  wire [31:0] _T_645; // @[Decode.scala 14:65]
  wire  _T_646; // @[Decode.scala 14:121]
  wire  _T_648; // @[Decode.scala 15:30]
  wire  _T_649; // @[Decode.scala 15:30]
  wire  _T_650; // @[Decode.scala 15:30]
  wire  _T_651; // @[Decode.scala 15:30]
  wire [3:0] id_ctrl_alu_fn; // @[Cat.scala 29:58]
  wire  _T_656; // @[Decode.scala 15:30]
  wire  _T_657; // @[Decode.scala 15:30]
  wire  _T_658; // @[Decode.scala 15:30]
  wire  _T_659; // @[Decode.scala 15:30]
  wire  _T_660; // @[Decode.scala 15:30]
  wire  _T_661; // @[Decode.scala 15:30]
  wire  _T_662; // @[Decode.scala 15:30]
  wire  _T_663; // @[Decode.scala 15:30]
  wire  _T_664; // @[Decode.scala 15:30]
  wire  _T_665; // @[Decode.scala 15:30]
  wire  _T_666; // @[Decode.scala 15:30]
  wire  _T_667; // @[Decode.scala 15:30]
  wire  _T_668; // @[Decode.scala 15:30]
  wire  _T_669; // @[Decode.scala 15:30]
  wire  _T_670; // @[Decode.scala 15:30]
  wire  _T_671; // @[Decode.scala 15:30]
  wire  _T_672; // @[Decode.scala 15:30]
  wire  _T_673; // @[Decode.scala 15:30]
  wire  _T_674; // @[Decode.scala 15:30]
  wire  _T_675; // @[Decode.scala 15:30]
  wire  _T_676; // @[Decode.scala 15:30]
  wire  _T_677; // @[Decode.scala 15:30]
  wire  _T_678; // @[Decode.scala 15:30]
  wire  _T_679; // @[Decode.scala 15:30]
  wire  _T_680; // @[Decode.scala 15:30]
  wire  _T_681; // @[Decode.scala 15:30]
  wire  _T_682; // @[Decode.scala 15:30]
  wire  _T_683; // @[Decode.scala 15:30]
  wire  _T_684; // @[Decode.scala 15:30]
  wire  _T_685; // @[Decode.scala 15:30]
  wire  _T_686; // @[Decode.scala 15:30]
  wire  _T_687; // @[Decode.scala 15:30]
  wire  _T_688; // @[Decode.scala 15:30]
  wire  _T_689; // @[Decode.scala 15:30]
  wire  _T_690; // @[Decode.scala 15:30]
  wire  _T_691; // @[Decode.scala 15:30]
  wire  id_ctrl_mem; // @[Decode.scala 15:30]
  wire  _T_694; // @[Decode.scala 14:121]
  wire [31:0] _T_695; // @[Decode.scala 14:65]
  wire  _T_696; // @[Decode.scala 14:121]
  wire [31:0] _T_697; // @[Decode.scala 14:65]
  wire  _T_698; // @[Decode.scala 14:121]
  wire  _T_700; // @[Decode.scala 15:30]
  wire  _T_701; // @[Decode.scala 15:30]
  wire [31:0] _T_702; // @[Decode.scala 14:65]
  wire  _T_703; // @[Decode.scala 14:121]
  wire [31:0] _T_704; // @[Decode.scala 14:65]
  wire  _T_705; // @[Decode.scala 14:121]
  wire  _T_707; // @[Decode.scala 15:30]
  wire [31:0] _T_708; // @[Decode.scala 14:65]
  wire  _T_709; // @[Decode.scala 14:121]
  wire [31:0] _T_710; // @[Decode.scala 14:65]
  wire  _T_711; // @[Decode.scala 14:121]
  wire [31:0] _T_712; // @[Decode.scala 14:65]
  wire  _T_713; // @[Decode.scala 14:121]
  wire  _T_715; // @[Decode.scala 15:30]
  wire  _T_716; // @[Decode.scala 15:30]
  wire  _T_717; // @[Decode.scala 15:30]
  wire [31:0] _T_718; // @[Decode.scala 14:65]
  wire  _T_719; // @[Decode.scala 14:121]
  wire [4:0] id_ctrl_mem_cmd; // @[Cat.scala 29:58]
  wire [31:0] _T_726; // @[Decode.scala 14:65]
  wire  _T_727; // @[Decode.scala 14:121]
  wire [31:0] _T_728; // @[Decode.scala 14:65]
  wire  _T_729; // @[Decode.scala 14:121]
  wire [31:0] _T_730; // @[Decode.scala 14:65]
  wire  id_ctrl_rfs3; // @[Decode.scala 14:121]
  wire  _T_733; // @[Decode.scala 15:30]
  wire  id_ctrl_rfs1; // @[Decode.scala 15:30]
  wire [31:0] _T_735; // @[Decode.scala 14:65]
  wire  _T_736; // @[Decode.scala 14:121]
  wire [31:0] _T_737; // @[Decode.scala 14:65]
  wire  _T_738; // @[Decode.scala 14:121]
  wire [31:0] _T_739; // @[Decode.scala 14:65]
  wire  _T_740; // @[Decode.scala 14:121]
  wire  _T_742; // @[Decode.scala 15:30]
  wire  _T_743; // @[Decode.scala 15:30]
  wire  id_ctrl_rfs2; // @[Decode.scala 15:30]
  wire [31:0] _T_746; // @[Decode.scala 14:65]
  wire  _T_747; // @[Decode.scala 14:121]
  wire  _T_749; // @[Decode.scala 14:121]
  wire  _T_751; // @[Decode.scala 15:30]
  wire  _T_752; // @[Decode.scala 15:30]
  wire  id_ctrl_wfd; // @[Decode.scala 15:30]
  wire [31:0] _T_754; // @[Decode.scala 14:65]
  wire  id_ctrl_div; // @[Decode.scala 14:121]
  wire  _T_758; // @[Decode.scala 14:121]
  wire  _T_760; // @[Decode.scala 14:121]
  wire [31:0] _T_761; // @[Decode.scala 14:65]
  wire  _T_762; // @[Decode.scala 14:121]
  wire [31:0] _T_763; // @[Decode.scala 14:65]
  wire  _T_764; // @[Decode.scala 14:121]
  wire [31:0] _T_765; // @[Decode.scala 14:65]
  wire  _T_766; // @[Decode.scala 14:121]
  wire [31:0] _T_767; // @[Decode.scala 14:65]
  wire  _T_768; // @[Decode.scala 14:121]
  wire [31:0] _T_769; // @[Decode.scala 14:65]
  wire  _T_770; // @[Decode.scala 14:121]
  wire  _T_772; // @[Decode.scala 15:30]
  wire  _T_773; // @[Decode.scala 15:30]
  wire  _T_774; // @[Decode.scala 15:30]
  wire  _T_775; // @[Decode.scala 15:30]
  wire  _T_776; // @[Decode.scala 15:30]
  wire  id_ctrl_wxd; // @[Decode.scala 15:30]
  wire [31:0] _T_778; // @[Decode.scala 14:65]
  wire  _T_779; // @[Decode.scala 14:121]
  wire [31:0] _T_781; // @[Decode.scala 14:65]
  wire  _T_782; // @[Decode.scala 14:121]
  wire [31:0] _T_784; // @[Decode.scala 14:65]
  wire  _T_785; // @[Decode.scala 14:121]
  wire [31:0] _T_786; // @[Decode.scala 14:65]
  wire  _T_787; // @[Decode.scala 14:121]
  wire [31:0] _T_788; // @[Decode.scala 14:65]
  wire  _T_789; // @[Decode.scala 14:121]
  wire  _T_791; // @[Decode.scala 15:30]
  wire  _T_792; // @[Decode.scala 15:30]
  wire  _T_793; // @[Decode.scala 15:30]
  wire  _T_794; // @[Decode.scala 15:30]
  wire [2:0] id_ctrl_csr; // @[Cat.scala 29:58]
  wire [31:0] _T_797; // @[Decode.scala 14:65]
  wire  id_ctrl_fence_i; // @[Decode.scala 14:121]
  wire  id_ctrl_fence; // @[Decode.scala 14:121]
  wire [31:0] _T_803; // @[Decode.scala 14:65]
  wire  id_ctrl_amo; // @[Decode.scala 14:121]
  wire [31:0] _T_806; // @[Decode.scala 14:65]
  wire  _T_807; // @[Decode.scala 14:121]
  wire [31:0] _T_808; // @[Decode.scala 14:65]
  wire  _T_809; // @[Decode.scala 14:121]
  wire [31:0] _T_810; // @[Decode.scala 14:65]
  wire  _T_811; // @[Decode.scala 14:121]
  wire  _T_813; // @[Decode.scala 15:30]
  wire  id_ctrl_dp; // @[Decode.scala 15:30]
  wire [4:0] id_raddr3; // @[RocketCore.scala 261:72]
  wire [4:0] id_raddr2; // @[RocketCore.scala 261:72]
  wire [4:0] id_raddr1; // @[RocketCore.scala 261:72]
  wire [4:0] id_waddr; // @[RocketCore.scala 261:72]
  reg  id_reg_fence; // @[RocketCore.scala 268:25]
  reg [31:0] _RAND_94;
  wire  _T_816; // @[RocketCore.scala 1021:45]
  wire [63:0] _T_821; // @[RocketCore.scala 1021:25]
  wire [63:0] _T_827; // @[RocketCore.scala 1021:25]
  wire  _T_894; // @[package.scala 15:47]
  wire  _T_895; // @[package.scala 15:47]
  wire  _T_896; // @[package.scala 15:47]
  wire  _T_897; // @[package.scala 64:59]
  wire  id_csr_en; // @[package.scala 64:59]
  wire  id_system_insn; // @[RocketCore.scala 278:36]
  wire  id_csr_ren; // @[RocketCore.scala 279:54]
  wire  _T_902; // @[RocketCore.scala 281:50]
  wire  id_sfence; // @[RocketCore.scala 281:31]
  wire  _T_903; // @[RocketCore.scala 282:32]
  wire  _T_905; // @[RocketCore.scala 282:64]
  wire  _T_906; // @[RocketCore.scala 282:79]
  wire  id_csr_flush; // @[RocketCore.scala 282:50]
  wire  _T_911; // @[RocketCore.scala 291:34]
  wire  _T_912; // @[RocketCore.scala 290:40]
  wire  _T_915; // @[RocketCore.scala 292:17]
  wire  _T_916; // @[RocketCore.scala 291:65]
  wire  _T_917; // @[RocketCore.scala 293:48]
  wire  _T_918; // @[RocketCore.scala 293:16]
  wire  _T_919; // @[RocketCore.scala 292:48]
  wire  _T_922; // @[RocketCore.scala 294:16]
  wire  _T_923; // @[RocketCore.scala 293:70]
  wire  _T_926; // @[RocketCore.scala 295:30]
  wire  _T_927; // @[RocketCore.scala 294:47]
  wire  _T_947; // @[RocketCore.scala 301:64]
  wire  _T_948; // @[RocketCore.scala 301:49]
  wire  _T_949; // @[RocketCore.scala 301:15]
  wire  _T_950; // @[RocketCore.scala 300:81]
  wire  _T_953; // @[RocketCore.scala 302:65]
  wire  _T_954; // @[RocketCore.scala 302:31]
  wire  id_illegal_insn; // @[RocketCore.scala 301:99]
  wire  id_amo_aq; // @[RocketCore.scala 304:29]
  wire  id_amo_rl; // @[RocketCore.scala 305:29]
  wire [3:0] id_fence_succ; // @[RocketCore.scala 307:33]
  wire  _T_955; // @[RocketCore.scala 308:52]
  wire  id_fence_next; // @[RocketCore.scala 308:37]
  wire  id_mem_busy; // @[RocketCore.scala 309:38]
  wire  _GEN_0; // @[RocketCore.scala 310:23]
  wire  _T_965; // @[RocketCore.scala 315:33]
  wire  _T_966; // @[RocketCore.scala 315:46]
  wire  _T_968; // @[RocketCore.scala 315:81]
  wire  _T_969; // @[RocketCore.scala 315:65]
  wire  id_do_fence; // @[RocketCore.scala 315:17]
  wire  _T_972; // @[RocketCore.scala 974:26]
  wire  _T_973; // @[RocketCore.scala 974:26]
  wire  _T_974; // @[RocketCore.scala 974:26]
  wire  _T_975; // @[RocketCore.scala 974:26]
  wire  _T_976; // @[RocketCore.scala 974:26]
  wire  _T_977; // @[RocketCore.scala 974:26]
  wire  id_xcpt; // @[RocketCore.scala 974:26]
  wire [1:0] _T_978; // @[Mux.scala 47:69]
  wire [3:0] _T_979; // @[Mux.scala 47:69]
  wire [3:0] _T_980; // @[Mux.scala 47:69]
  wire [3:0] _T_981; // @[Mux.scala 47:69]
  wire [3:0] _T_982; // @[Mux.scala 47:69]
  wire [3:0] _T_983; // @[Mux.scala 47:69]
  wire [4:0] ex_waddr; // @[RocketCore.scala 351:29]
  wire [4:0] mem_waddr; // @[RocketCore.scala 352:31]
  wire [4:0] wb_waddr; // @[RocketCore.scala 353:29]
  wire  _T_997; // @[RocketCore.scala 356:19]
  wire  _T_998; // @[RocketCore.scala 357:20]
  wire  _T_1000; // @[RocketCore.scala 357:36]
  wire  id_bypass_src_0_0; // @[RocketCore.scala 359:82]
  wire  _T_1003; // @[RocketCore.scala 359:82]
  wire  id_bypass_src_0_1; // @[RocketCore.scala 359:74]
  wire  _T_1004; // @[RocketCore.scala 359:82]
  wire  id_bypass_src_0_2; // @[RocketCore.scala 359:74]
  wire  id_bypass_src_0_3; // @[RocketCore.scala 359:74]
  wire  id_bypass_src_1_0; // @[RocketCore.scala 359:82]
  wire  _T_1007; // @[RocketCore.scala 359:82]
  wire  id_bypass_src_1_1; // @[RocketCore.scala 359:74]
  wire  _T_1008; // @[RocketCore.scala 359:82]
  wire  id_bypass_src_1_2; // @[RocketCore.scala 359:74]
  wire  id_bypass_src_1_3; // @[RocketCore.scala 359:74]
  reg  ex_reg_rs_bypass_0; // @[RocketCore.scala 363:29]
  reg [31:0] _RAND_95;
  reg  ex_reg_rs_bypass_1; // @[RocketCore.scala 363:29]
  reg [31:0] _RAND_96;
  reg [1:0] ex_reg_rs_lsb_0; // @[RocketCore.scala 364:26]
  reg [31:0] _RAND_97;
  reg [1:0] ex_reg_rs_lsb_1; // @[RocketCore.scala 364:26]
  reg [31:0] _RAND_98;
  reg [61:0] ex_reg_rs_msb_0; // @[RocketCore.scala 365:26]
  reg [63:0] _RAND_99;
  reg [61:0] ex_reg_rs_msb_1; // @[RocketCore.scala 365:26]
  reg [63:0] _RAND_100;
  wire  _T_1010; // @[package.scala 32:86]
  wire [63:0] _T_1011; // @[package.scala 32:76]
  wire  _T_1012; // @[package.scala 32:86]
  wire [63:0] _T_1013; // @[package.scala 32:76]
  wire  _T_1014; // @[package.scala 32:86]
  wire [63:0] _T_1015; // @[package.scala 32:76]
  wire [63:0] _T_1016; // @[Cat.scala 29:58]
  wire  _T_1017; // @[package.scala 32:86]
  wire [63:0] _T_1018; // @[package.scala 32:76]
  wire  _T_1019; // @[package.scala 32:86]
  wire [63:0] _T_1020; // @[package.scala 32:76]
  wire  _T_1021; // @[package.scala 32:86]
  wire [63:0] _T_1022; // @[package.scala 32:76]
  wire [63:0] _T_1023; // @[Cat.scala 29:58]
  wire [63:0] ex_rs_1; // @[RocketCore.scala 367:14]
  wire  _T_1024; // @[RocketCore.scala 1036:24]
  wire  _T_1026; // @[RocketCore.scala 1036:53]
  wire  _T_1027; // @[RocketCore.scala 1036:19]
  wire  _T_1028; // @[RocketCore.scala 1037:26]
  wire [10:0] _T_1030; // @[RocketCore.scala 1037:49]
  wire  _T_1032; // @[RocketCore.scala 1038:26]
  wire  _T_1033; // @[RocketCore.scala 1038:43]
  wire  _T_1034; // @[RocketCore.scala 1038:36]
  wire [7:0] _T_1036; // @[RocketCore.scala 1038:73]
  wire  _T_1040; // @[RocketCore.scala 1039:33]
  wire  _T_1041; // @[RocketCore.scala 1040:23]
  wire  _T_1043; // @[RocketCore.scala 1040:44]
  wire  _T_1044; // @[RocketCore.scala 1041:23]
  wire  _T_1046; // @[RocketCore.scala 1041:43]
  wire  _T_1047; // @[RocketCore.scala 1041:18]
  wire  _T_1048; // @[RocketCore.scala 1040:18]
  wire [5:0] _T_1054; // @[RocketCore.scala 1042:20]
  wire  _T_1056; // @[RocketCore.scala 1044:24]
  wire  _T_1058; // @[RocketCore.scala 1044:34]
  wire [3:0] _T_1063; // @[RocketCore.scala 1045:19]
  wire [3:0] _T_1064; // @[RocketCore.scala 1044:19]
  wire [3:0] _T_1065; // @[RocketCore.scala 1043:19]
  wire  _T_1068; // @[RocketCore.scala 1047:22]
  wire  _T_1072; // @[RocketCore.scala 1048:17]
  wire  _T_1073; // @[RocketCore.scala 1047:17]
  wire  _T_1074; // @[RocketCore.scala 1046:17]
  wire  _T_1077; // @[Cat.scala 29:58]
  wire [7:0] _T_1078; // @[Cat.scala 29:58]
  wire [10:0] _T_1080; // @[Cat.scala 29:58]
  wire  _T_1081; // @[Cat.scala 29:58]
  wire [31:0] ex_imm; // @[RocketCore.scala 1050:53]
  wire [63:0] _T_1085; // @[RocketCore.scala 370:24]
  wire  _T_1087; // @[Mux.scala 80:60]
  wire [63:0] _T_1088; // @[Mux.scala 80:57]
  wire  _T_1089; // @[Mux.scala 80:60]
  wire [63:0] _T_1090; // @[RocketCore.scala 373:24]
  wire [3:0] _T_1091; // @[RocketCore.scala 375:19]
  wire  _T_1092; // @[Mux.scala 80:60]
  wire [63:0] _T_1093; // @[Mux.scala 80:57]
  wire  _T_1094; // @[Mux.scala 80:60]
  wire [63:0] _T_1095; // @[Mux.scala 80:57]
  wire  _T_1096; // @[Mux.scala 80:60]
  wire  _T_1763; // @[RocketCore.scala 776:40]
  wire  _T_1764; // @[RocketCore.scala 776:71]
  wire  _T_1568; // @[RocketCore.scala 706:55]
  wire  _T_1569; // @[RocketCore.scala 706:42]
  wire  _T_1616; // @[RocketCore.scala 726:70]
  wire  _T_1617; // @[RocketCore.scala 983:27]
  wire  _T_1570; // @[RocketCore.scala 707:55]
  wire  _T_1571; // @[RocketCore.scala 707:42]
  wire  _T_1618; // @[RocketCore.scala 726:70]
  wire  _T_1619; // @[RocketCore.scala 983:27]
  wire  _T_1622; // @[RocketCore.scala 983:50]
  wire  _T_1572; // @[RocketCore.scala 708:55]
  wire  _T_1573; // @[RocketCore.scala 708:42]
  wire  _T_1620; // @[RocketCore.scala 726:70]
  wire  _T_1621; // @[RocketCore.scala 983:27]
  wire  _T_1623; // @[RocketCore.scala 983:50]
  wire  data_hazard_ex; // @[RocketCore.scala 726:36]
  wire  _T_1609; // @[RocketCore.scala 725:38]
  wire  _T_1610; // @[RocketCore.scala 725:48]
  wire  _T_1611; // @[RocketCore.scala 725:64]
  wire  _T_1613; // @[RocketCore.scala 725:94]
  wire  ex_cannot_bypass; // @[RocketCore.scala 725:109]
  wire  _T_1635; // @[RocketCore.scala 728:54]
  wire  _T_1625; // @[RocketCore.scala 983:27]
  wire  _T_1627; // @[RocketCore.scala 983:27]
  wire  _T_1632; // @[RocketCore.scala 983:50]
  wire  _T_1628; // @[RocketCore.scala 727:76]
  wire  _T_1629; // @[RocketCore.scala 983:27]
  wire  _T_1633; // @[RocketCore.scala 983:50]
  wire  _T_1631; // @[RocketCore.scala 983:27]
  wire  _T_1634; // @[RocketCore.scala 983:50]
  wire  fp_data_hazard_ex; // @[RocketCore.scala 727:39]
  wire  _T_1636; // @[RocketCore.scala 728:74]
  wire  id_ex_hazard; // @[RocketCore.scala 728:35]
  wire  _T_1643; // @[RocketCore.scala 735:72]
  wire  _T_1644; // @[RocketCore.scala 983:27]
  wire  _T_1645; // @[RocketCore.scala 735:72]
  wire  _T_1646; // @[RocketCore.scala 983:27]
  wire  _T_1649; // @[RocketCore.scala 983:50]
  wire  _T_1647; // @[RocketCore.scala 735:72]
  wire  _T_1648; // @[RocketCore.scala 983:27]
  wire  _T_1650; // @[RocketCore.scala 983:50]
  wire  data_hazard_mem; // @[RocketCore.scala 735:38]
  wire  _T_1637; // @[RocketCore.scala 734:40]
  wire  _T_1638; // @[RocketCore.scala 734:66]
  wire  _T_1639; // @[RocketCore.scala 734:50]
  wire  _T_1641; // @[RocketCore.scala 734:100]
  wire  mem_cannot_bypass; // @[RocketCore.scala 734:116]
  wire  _T_1662; // @[RocketCore.scala 737:57]
  wire  _T_1652; // @[RocketCore.scala 983:27]
  wire  _T_1654; // @[RocketCore.scala 983:27]
  wire  _T_1659; // @[RocketCore.scala 983:50]
  wire  _T_1655; // @[RocketCore.scala 736:78]
  wire  _T_1656; // @[RocketCore.scala 983:27]
  wire  _T_1660; // @[RocketCore.scala 983:50]
  wire  _T_1658; // @[RocketCore.scala 983:27]
  wire  _T_1661; // @[RocketCore.scala 983:50]
  wire  fp_data_hazard_mem; // @[RocketCore.scala 736:41]
  wire  _T_1663; // @[RocketCore.scala 737:78]
  wire  id_mem_hazard; // @[RocketCore.scala 737:37]
  wire  _T_1733; // @[RocketCore.scala 764:18]
  wire  _T_1666; // @[RocketCore.scala 741:70]
  wire  _T_1667; // @[RocketCore.scala 983:27]
  wire  _T_1668; // @[RocketCore.scala 741:70]
  wire  _T_1669; // @[RocketCore.scala 983:27]
  wire  _T_1672; // @[RocketCore.scala 983:50]
  wire  _T_1670; // @[RocketCore.scala 741:70]
  wire  _T_1671; // @[RocketCore.scala 983:27]
  wire  _T_1673; // @[RocketCore.scala 983:50]
  wire  data_hazard_wb; // @[RocketCore.scala 741:36]
  wire  wb_dcache_miss; // @[RocketCore.scala 483:36]
  wire  wb_set_sboard; // @[RocketCore.scala 628:35]
  wire  _T_1685; // @[RocketCore.scala 743:54]
  wire  _T_1675; // @[RocketCore.scala 983:27]
  wire  _T_1677; // @[RocketCore.scala 983:27]
  wire  _T_1682; // @[RocketCore.scala 983:50]
  wire  _T_1678; // @[RocketCore.scala 742:76]
  wire  _T_1679; // @[RocketCore.scala 983:27]
  wire  _T_1683; // @[RocketCore.scala 983:50]
  wire  _T_1681; // @[RocketCore.scala 983:27]
  wire  _T_1684; // @[RocketCore.scala 983:50]
  wire  fp_data_hazard_wb; // @[RocketCore.scala 742:39]
  wire  _T_1686; // @[RocketCore.scala 743:71]
  wire  id_wb_hazard; // @[RocketCore.scala 743:35]
  wire  _T_1734; // @[RocketCore.scala 764:35]
  reg [31:0] _T_1574; // @[RocketCore.scala 1000:25]
  reg [31:0] _RAND_101;
  wire [31:0] _T_1576; // @[RocketCore.scala 1001:40]
  wire [31:0] _T_1582; // @[RocketCore.scala 997:35]
  wire  dmem_resp_valid; // @[RocketCore.scala 638:44]
  wire  dmem_resp_replay; // @[RocketCore.scala 639:42]
  wire  dmem_resp_xpu; // @[RocketCore.scala 635:23]
  wire  _T_1511; // @[RocketCore.scala 654:26]
  wire  _T_1510; // @[Decoupled.scala 40:37]
  wire  ll_wen; // @[RocketCore.scala 654:44]
  wire [4:0] dmem_resp_waddr; // @[RocketCore.scala 637:46]
  wire [4:0] ll_waddr; // @[RocketCore.scala 654:44]
  wire  _T_1584; // @[RocketCore.scala 718:70]
  wire  _T_1585; // @[RocketCore.scala 718:58]
  wire  _T_1587; // @[RocketCore.scala 721:77]
  wire  _T_1588; // @[RocketCore.scala 983:27]
  wire [31:0] _T_1589; // @[RocketCore.scala 997:35]
  wire  _T_1591; // @[RocketCore.scala 718:70]
  wire  _T_1592; // @[RocketCore.scala 718:58]
  wire  _T_1594; // @[RocketCore.scala 721:77]
  wire  _T_1595; // @[RocketCore.scala 983:27]
  wire  _T_1603; // @[RocketCore.scala 983:50]
  wire [31:0] _T_1596; // @[RocketCore.scala 997:35]
  wire  _T_1598; // @[RocketCore.scala 718:70]
  wire  _T_1599; // @[RocketCore.scala 718:58]
  wire  _T_1601; // @[RocketCore.scala 721:77]
  wire  _T_1602; // @[RocketCore.scala 983:27]
  wire  id_sboard_hazard; // @[RocketCore.scala 983:50]
  wire  _T_1735; // @[RocketCore.scala 764:51]
  wire  _T_1736; // @[RocketCore.scala 765:40]
  wire  _T_1737; // @[RocketCore.scala 765:57]
  wire  _T_1738; // @[RocketCore.scala 765:23]
  wire  _T_1739; // @[RocketCore.scala 764:71]
  wire  _T_1740; // @[RocketCore.scala 766:15]
  wire  _T_1742; // @[RocketCore.scala 766:42]
  wire  _T_1743; // @[RocketCore.scala 765:74]
  reg [31:0] _T_1687; // @[RocketCore.scala 1000:25]
  reg [31:0] _RAND_102;
  wire [31:0] _T_1706; // @[RocketCore.scala 997:35]
  wire  _T_1708; // @[RocketCore.scala 983:27]
  wire [31:0] _T_1709; // @[RocketCore.scala 997:35]
  wire  _T_1711; // @[RocketCore.scala 983:27]
  wire  _T_1718; // @[RocketCore.scala 983:50]
  wire [31:0] _T_1712; // @[RocketCore.scala 997:35]
  wire  _T_1714; // @[RocketCore.scala 983:27]
  wire  _T_1719; // @[RocketCore.scala 983:50]
  wire [31:0] _T_1715; // @[RocketCore.scala 997:35]
  wire  _T_1717; // @[RocketCore.scala 983:27]
  wire  id_stall_fpu; // @[RocketCore.scala 983:50]
  wire  _T_1744; // @[RocketCore.scala 767:16]
  wire  _T_1745; // @[RocketCore.scala 766:62]
  reg  blocked; // @[RocketCore.scala 756:22]
  reg [31:0] _RAND_103;
  wire  dcache_blocked; // @[RocketCore.scala 758:13]
  wire  _T_1746; // @[RocketCore.scala 768:17]
  wire  _T_1747; // @[RocketCore.scala 767:32]
  wire  wb_wxd; // @[RocketCore.scala 627:29]
  wire  _T_1751; // @[RocketCore.scala 770:62]
  wire  _T_1752; // @[RocketCore.scala 770:40]
  wire  _T_1754; // @[RocketCore.scala 770:75]
  wire  _T_1755; // @[RocketCore.scala 770:17]
  wire  _T_1756; // @[RocketCore.scala 769:34]
  wire  _T_1759; // @[RocketCore.scala 771:15]
  wire  _T_1760; // @[RocketCore.scala 772:17]
  wire  ctrl_stalld; // @[RocketCore.scala 773:22]
  wire  _T_1765; // @[RocketCore.scala 776:89]
  wire  ctrl_killd; // @[RocketCore.scala 776:104]
  wire  _T_1102; // @[RocketCore.scala 416:29]
  wire  _T_1112; // @[RocketCore.scala 426:42]
  wire  _T_1113; // @[RocketCore.scala 426:25]
  wire  _GEN_1; // @[RocketCore.scala 426:49]
  wire  _GEN_2; // @[RocketCore.scala 427:26]
  wire [1:0] _T_1114; // @[RocketCore.scala 433:22]
  wire  _T_1115; // @[RocketCore.scala 433:29]
  wire  _GEN_5; // @[RocketCore.scala 433:34]
  wire [1:0] _T_1116; // @[RocketCore.scala 438:40]
  wire  _T_1117; // @[RocketCore.scala 438:47]
  wire  _T_1118; // @[RocketCore.scala 438:28]
  wire  _GEN_9; // @[RocketCore.scala 428:20]
  wire  _T_1119; // @[RocketCore.scala 443:42]
  wire  _T_1122; // @[package.scala 15:47]
  wire  _T_1123; // @[package.scala 64:59]
  wire [1:0] _T_1126; // @[Cat.scala 29:58]
  wire  _T_1127; // @[RocketCore.scala 456:48]
  wire  _T_1128; // @[RocketCore.scala 456:48]
  wire  do_bypass; // @[RocketCore.scala 456:48]
  wire  _T_1132; // @[RocketCore.scala 460:23]
  wire  _T_1513; // @[RocketCore.scala 662:31]
  wire  wb_valid; // @[RocketCore.scala 662:45]
  wire  wb_wen; // @[RocketCore.scala 663:25]
  wire  rf_wen; // @[RocketCore.scala 664:23]
  wire [4:0] rf_waddr; // @[RocketCore.scala 665:21]
  wire  _T_1521; // @[RocketCore.scala 1026:16]
  wire  _T_1525; // @[RocketCore.scala 1029:20]
  wire  _T_1515; // @[RocketCore.scala 666:38]
  wire [63:0] ll_wdata;
  wire  _T_1517; // @[RocketCore.scala 668:34]
  wire [63:0] _T_1519; // @[RocketCore.scala 668:21]
  wire [63:0] _T_1520; // @[RocketCore.scala 667:21]
  wire [63:0] rf_wdata; // @[RocketCore.scala 666:21]
  wire [63:0] _GEN_226; // @[RocketCore.scala 1029:31]
  wire [63:0] _GEN_233; // @[RocketCore.scala 1026:29]
  wire [63:0] id_rs_0; // @[RocketCore.scala 671:17]
  wire  _T_1135; // @[RocketCore.scala 456:48]
  wire  _T_1136; // @[RocketCore.scala 456:48]
  wire  do_bypass_1; // @[RocketCore.scala 456:48]
  wire  _T_1140; // @[RocketCore.scala 460:23]
  wire  _T_1526; // @[RocketCore.scala 1029:20]
  wire [63:0] _GEN_227; // @[RocketCore.scala 1029:31]
  wire [63:0] _GEN_234; // @[RocketCore.scala 1026:29]
  wire [63:0] id_rs_1; // @[RocketCore.scala 671:17]
  wire [31:0] inst; // @[RocketCore.scala 466:21]
  wire  _T_1664; // @[RocketCore.scala 738:32]
  wire  id_load_use; // @[RocketCore.scala 738:51]
  wire  _T_1147; // @[RocketCore.scala 472:21]
  wire  _T_1148; // @[RocketCore.scala 472:41]
  wire  _T_1152; // @[RocketCore.scala 484:42]
  wire  _T_1154; // @[RocketCore.scala 485:42]
  wire  replay_ex_structural; // @[RocketCore.scala 484:64]
  wire  replay_ex_load_use; // @[RocketCore.scala 486:43]
  wire  _T_1155; // @[RocketCore.scala 487:75]
  wire  _T_1156; // @[RocketCore.scala 487:50]
  wire  replay_ex; // @[RocketCore.scala 487:33]
  wire  _T_1157; // @[RocketCore.scala 488:35]
  wire  ctrl_killx; // @[RocketCore.scala 488:48]
  wire  _T_1159; // @[RocketCore.scala 490:40]
  wire  _T_1160; // @[RocketCore.scala 490:69]
  wire  ex_slow_bypass; // @[RocketCore.scala 490:50]
  wire  _T_1162; // @[RocketCore.scala 491:67]
  wire  ex_sfence; // @[RocketCore.scala 491:48]
  wire  ex_xcpt; // @[RocketCore.scala 494:28]
  wire  _T_1173; // @[RocketCore.scala 500:36]
  wire  mem_pc_valid; // @[RocketCore.scala 500:54]
  wire  _T_1326; // @[RocketCore.scala 509:56]
  wire  mem_npc_misaligned; // @[RocketCore.scala 509:70]
  wire  _T_1329; // @[RocketCore.scala 510:59]
  wire  _T_1330; // @[RocketCore.scala 510:41]
  wire [63:0] mem_int_wdata; // @[RocketCore.scala 510:119]
  wire  _T_1333; // @[RocketCore.scala 511:33]
  wire  mem_cfi; // @[RocketCore.scala 511:50]
  wire  _T_1335; // @[RocketCore.scala 512:57]
  wire  mem_cfi_taken; // @[RocketCore.scala 512:74]
  wire  _T_1347; // @[RocketCore.scala 524:23]
  wire  _T_1348; // @[Consts.scala 82:31]
  wire  _T_1349; // @[Consts.scala 82:48]
  wire  _T_1350; // @[Consts.scala 82:41]
  wire  _T_1352; // @[Consts.scala 82:58]
  wire  _T_1353; // @[package.scala 15:47]
  wire  _T_1354; // @[package.scala 15:47]
  wire  _T_1355; // @[package.scala 15:47]
  wire  _T_1356; // @[package.scala 15:47]
  wire  _T_1357; // @[package.scala 64:59]
  wire  _T_1358; // @[package.scala 64:59]
  wire  _T_1359; // @[package.scala 64:59]
  wire  _T_1360; // @[package.scala 15:47]
  wire  _T_1361; // @[package.scala 15:47]
  wire  _T_1362; // @[package.scala 15:47]
  wire  _T_1363; // @[package.scala 15:47]
  wire  _T_1364; // @[package.scala 15:47]
  wire  _T_1365; // @[package.scala 64:59]
  wire  _T_1366; // @[package.scala 64:59]
  wire  _T_1367; // @[package.scala 64:59]
  wire  _T_1368; // @[package.scala 64:59]
  wire  _T_1369; // @[Consts.scala 80:44]
  wire  _T_1370; // @[Consts.scala 82:75]
  wire  _T_1371; // @[RocketCore.scala 531:33]
  wire  _T_1372; // @[Consts.scala 83:32]
  wire  _T_1373; // @[Consts.scala 83:49]
  wire  _T_1374; // @[Consts.scala 83:42]
  wire  _T_1376; // @[Consts.scala 83:59]
  wire  _T_1394; // @[Consts.scala 83:76]
  wire  _T_1395; // @[RocketCore.scala 532:34]
  wire [63:0] _T_1396; // @[RocketCore.scala 544:25]
  wire  _T_1398; // @[RocketCore.scala 547:56]
  wire  _T_1399; // @[RocketCore.scala 547:24]
  wire  _T_1401; // @[AMOALU.scala 26:19]
  wire [63:0] _T_1405; // @[Cat.scala 29:58]
  wire  _T_1406; // @[AMOALU.scala 26:19]
  wire [63:0] _T_1409; // @[Cat.scala 29:58]
  wire  _T_1410; // @[AMOALU.scala 26:19]
  wire [63:0] _T_1412; // @[Cat.scala 29:58]
  wire  _T_1416; // @[RocketCore.scala 551:24]
  wire  _GEN_77; // @[RocketCore.scala 551:48]
  wire  _GEN_78; // @[RocketCore.scala 551:48]
  wire  _T_1417; // @[RocketCore.scala 558:38]
  wire  _T_1418; // @[RocketCore.scala 558:75]
  wire  mem_breakpoint; // @[RocketCore.scala 558:57]
  wire  _T_1419; // @[RocketCore.scala 559:44]
  wire  _T_1420; // @[RocketCore.scala 559:82]
  wire  mem_debug_breakpoint; // @[RocketCore.scala 559:64]
  wire  mem_ldst_xcpt; // @[RocketCore.scala 974:26]
  wire [3:0] mem_ldst_cause; // @[Mux.scala 47:69]
  wire  _T_1421; // @[RocketCore.scala 565:29]
  wire  _T_1422; // @[RocketCore.scala 566:20]
  wire  _T_1423; // @[RocketCore.scala 567:20]
  wire  _T_1424; // @[RocketCore.scala 974:26]
  wire  mem_xcpt; // @[RocketCore.scala 974:26]
  wire [3:0] _T_1425; // @[Mux.scala 47:69]
  wire  dcache_kill_mem; // @[RocketCore.scala 576:55]
  wire  _T_1439; // @[RocketCore.scala 577:36]
  wire  fpu_kill_mem; // @[RocketCore.scala 577:51]
  wire  _T_1440; // @[RocketCore.scala 578:37]
  wire  replay_mem; // @[RocketCore.scala 578:55]
  wire  _T_1441; // @[RocketCore.scala 579:38]
  wire  _T_1442; // @[RocketCore.scala 579:52]
  wire  killm_common; // @[RocketCore.scala 579:68]
  reg  _T_1445; // @[RocketCore.scala 580:37]
  reg [31:0] _RAND_104;
  wire  _T_1447; // @[RocketCore.scala 581:33]
  wire  ctrl_killm; // @[RocketCore.scala 581:45]
  wire  _T_1456; // @[RocketCore.scala 592:25]
  wire  _T_1457; // @[RocketCore.scala 592:40]
  wire [2:0] _T_1482; // @[Mux.scala 47:69]
  wire [3:0] _T_1483; // @[Mux.scala 47:69]
  wire [3:0] _T_1484; // @[Mux.scala 47:69]
  wire [3:0] _T_1485; // @[Mux.scala 47:69]
  wire [3:0] _T_1486; // @[Mux.scala 47:69]
  wire [63:0] wb_cause; // @[Mux.scala 47:69]
  wire  _T_1487; // @[RocketCore.scala 978:38]
  wire  _T_1489; // @[RocketCore.scala 978:38]
  wire  _T_1491; // @[RocketCore.scala 978:38]
  wire  _T_1493; // @[RocketCore.scala 978:38]
  wire  _T_1495; // @[RocketCore.scala 978:38]
  wire  _T_1497; // @[RocketCore.scala 978:38]
  wire  _T_1529; // @[RocketCore.scala 679:73]
  wire [15:0] _T_1531; // @[RocketCore.scala 679:50]
  wire  _T_1535; // @[package.scala 15:47]
  wire  _T_1536; // @[package.scala 15:47]
  wire  _T_1541; // @[package.scala 15:47]
  wire  _T_1544; // @[package.scala 15:47]
  wire  _T_1545; // @[package.scala 64:59]
  wire  _T_1546; // @[package.scala 64:59]
  wire  _T_1547; // @[package.scala 64:59]
  wire  _T_1548; // @[package.scala 64:59]
  wire  _T_1549; // @[package.scala 64:59]
  wire  _T_1550; // @[package.scala 64:59]
  wire  _T_1551; // @[package.scala 64:59]
  wire  _T_1552; // @[package.scala 64:59]
  wire  _T_1553; // @[package.scala 64:59]
  wire  tval_valid; // @[RocketCore.scala 688:28]
  wire [24:0] a_1; // @[RocketCore.scala 988:23]
  wire  _T_1555; // @[RocketCore.scala 989:21]
  wire  _T_1556; // @[RocketCore.scala 989:34]
  wire  _T_1557; // @[RocketCore.scala 989:29]
  wire  msb_1; // @[RocketCore.scala 989:18]
  wire [39:0] _T_1562; // @[Cat.scala 29:58]
  wire [2:0] _T_1565; // @[CSR.scala 131:15]
  wire [31:0] _T_1577; // @[RocketCore.scala 1004:62]
  wire [31:0] _T_1578; // @[RocketCore.scala 1004:49]
  wire [31:0] _T_1580; // @[RocketCore.scala 996:62]
  wire  _T_1604; // @[RocketCore.scala 722:28]
  wire [31:0] _T_1605; // @[RocketCore.scala 1004:62]
  wire [31:0] _T_1606; // @[RocketCore.scala 1004:49]
  wire [31:0] _T_1607; // @[RocketCore.scala 995:60]
  wire  _T_1608; // @[RocketCore.scala 1007:17]
  wire  _T_1688; // @[RocketCore.scala 747:35]
  wire  _T_1689; // @[RocketCore.scala 747:50]
  wire  _T_1690; // @[RocketCore.scala 747:72]
  wire [31:0] _T_1692; // @[RocketCore.scala 1004:49]
  wire [31:0] _T_1693; // @[RocketCore.scala 995:60]
  wire  _T_1695; // @[RocketCore.scala 748:38]
  wire [31:0] _T_1696; // @[RocketCore.scala 1004:62]
  wire [31:0] _T_1697; // @[RocketCore.scala 1004:49]
  wire [31:0] _T_1699; // @[RocketCore.scala 996:62]
  wire  _T_1700; // @[RocketCore.scala 1007:17]
  wire [31:0] _T_1701; // @[RocketCore.scala 1004:62]
  wire [31:0] _T_1702; // @[RocketCore.scala 1004:49]
  wire [31:0] _T_1704; // @[RocketCore.scala 996:62]
  wire  _T_1705; // @[RocketCore.scala 1007:17]
  wire  _T_1723; // @[RocketCore.scala 757:60]
  wire  _T_1724; // @[RocketCore.scala 757:95]
  wire  _T_1725; // @[RocketCore.scala 757:116]
  wire  _T_1768; // @[RocketCore.scala 781:17]
  wire [39:0] _T_1769; // @[RocketCore.scala 782:8]
  wire  _T_1771; // @[RocketCore.scala 784:40]
  wire  _T_1774; // @[RocketCore.scala 786:43]
  wire  _T_1782; // @[RocketCore.scala 798:45]
  wire  _T_1783; // @[RocketCore.scala 798:60]
  wire  _T_1785; // @[RocketCore.scala 798:90]
  wire  _T_1787; // @[RocketCore.scala 801:23]
  wire  _T_1789; // @[RocketCore.scala 801:41]
  wire [4:0] _T_1792; // @[RocketCore.scala 802:62]
  wire  _T_1793; // @[RocketCore.scala 802:62]
  wire  _T_1794; // @[RocketCore.scala 802:23]
  wire [1:0] _T_1797; // @[RocketCore.scala 802:8]
  wire [1:0] _T_1799; // @[RocketCore.scala 806:74]
  wire [39:0] _GEN_250; // @[RocketCore.scala 806:69]
  wire [39:0] _T_1801; // @[RocketCore.scala 806:69]
  wire [38:0] _T_1803; // @[RocketCore.scala 807:66]
  wire [5:0] ex_dcache_tag; // @[Cat.scala 29:58]
  wire [24:0] a_2; // @[RocketCore.scala 988:23]
  wire  _T_1815; // @[RocketCore.scala 989:21]
  wire  _T_1816; // @[RocketCore.scala 989:34]
  wire  _T_1817; // @[RocketCore.scala 989:29]
  wire  msb_2; // @[RocketCore.scala 989:18]
  wire  _T_1824; // @[RocketCore.scala 839:35]
  wire  _T_1845; // @[RocketCore.scala 852:62]
  wire  _T_1846; // @[RocketCore.scala 852:68]
  wire  unpause; // @[RocketCore.scala 852:92]
  wire  _T_1849; // @[RocketCore.scala 871:33]
  wire  coreMonitorBundle_valid; // @[RocketCore.scala 888:52]
  wire [39:0] _T_1858; // @[RocketCore.scala 889:48]
  wire [23:0] _T_1861; // @[Bitwise.scala 72:12]
  wire [63:0] coreMonitorBundle_pc; // @[Cat.scala 29:58]
  wire  coreMonitorBundle_wrenx; // @[RocketCore.scala 890:37]
  reg [63:0] _T_1866; // @[RocketCore.scala 895:43]
  reg [63:0] _RAND_105;
  reg [63:0] coreMonitorBundle_rd0val; // @[RocketCore.scala 895:34]
  reg [63:0] _RAND_106;
  reg [63:0] _T_1869; // @[RocketCore.scala 897:43]
  reg [63:0] _RAND_107;
  reg [63:0] coreMonitorBundle_rd1val; // @[RocketCore.scala 897:34]
  reg [63:0] _RAND_108;
  wire  _T_1871; // @[RocketCore.scala 933:26]
  wire [4:0] _T_1872; // @[RocketCore.scala 933:13]
  wire [63:0] _T_1873; // @[RocketCore.scala 934:13]
  wire  _T_1874; // @[RocketCore.scala 936:27]
  wire [4:0] _T_1875; // @[RocketCore.scala 936:13]
  wire [63:0] _T_1877; // @[RocketCore.scala 937:13]
  wire  _T_1878; // @[RocketCore.scala 938:27]
  wire [4:0] _T_1879; // @[RocketCore.scala 938:13]
  wire [63:0] _T_1881; // @[RocketCore.scala 939:13]
  wire [31:0] coreMonitorBundle_inst; // @[RocketCore.scala 882:31 RocketCore.scala 898:26]
  reg [19:0] Rocket_state; // @[Register tracking Rocket state]
  reg [31:0] _RAND_109;
  reg  Rocket_cov [0:1048575]; // @[Coverage map for Rocket]
  reg [31:0] _RAND_110;
  wire  Rocket_cov_read_data; // @[Coverage map for Rocket]
  wire [19:0] Rocket_cov_read_addr; // @[Coverage map for Rocket]
  wire  Rocket_cov_write_data; // @[Coverage map for Rocket]
  wire [19:0] Rocket_cov_write_addr; // @[Coverage map for Rocket]
  wire  Rocket_cov_write_mask; // @[Coverage map for Rocket]
  wire  Rocket_cov_write_en; // @[Coverage map for Rocket]
  reg [29:0] Rocket_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_111;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire [16:0] mem_reg_slow_bypass_shl;
  wire [19:0] mem_reg_slow_bypass_pad;
  wire [1:0] ex_ctrl_sel_alu1_shl;
  wire [19:0] ex_ctrl_sel_alu1_pad;
  wire [2:0] ex_ctrl_wxd_shl;
  wire [19:0] ex_ctrl_wxd_pad;
  wire [18:0] wb_ctrl_rxs2_shl;
  wire [19:0] wb_ctrl_rxs2_pad;
  wire [16:0] mem_reg_store_shl;
  wire [19:0] mem_reg_store_pad;
  wire [6:0] wb_reg_valid_shl;
  wire [19:0] wb_reg_valid_pad;
  wire [2:0] mem_ctrl_jal_shl;
  wire [19:0] mem_ctrl_jal_pad;
  wire [16:0] mem_br_taken_shl;
  wire [19:0] mem_br_taken_pad;
  wire [13:0] ex_ctrl_jalr_shl;
  wire [19:0] ex_ctrl_jalr_pad;
  wire [11:0] wb_ctrl_rfs2_shl;
  wire [19:0] wb_ctrl_rfs2_pad;
  wire [9:0] ex_ctrl_sel_imm_shl;
  wire [19:0] ex_ctrl_sel_imm_pad;
  wire  mem_ctrl_mem_shl;
  wire [19:0] mem_ctrl_mem_pad;
  wire [6:0] wb_reg_xcpt_shl;
  wire [19:0] wb_reg_xcpt_pad;
  wire [11:0] ex_reg_xcpt_interrupt_shl;
  wire [19:0] ex_reg_xcpt_interrupt_pad;
  wire [9:0] mem_ctrl_branch_shl;
  wire [19:0] mem_ctrl_branch_pad;
  wire  ex_ctrl_fp_shl;
  wire [19:0] ex_ctrl_fp_pad;
  wire [9:0] ex_reg_mem_size_shl;
  wire [19:0] ex_reg_mem_size_pad;
  wire [1:0] mem_ctrl_wfd_shl;
  wire [19:0] mem_ctrl_wfd_pad;
  wire [18:0] mem_reg_load_shl;
  wire [19:0] mem_reg_load_pad;
  wire [18:0] mem_reg_flush_pipe_shl;
  wire [19:0] mem_reg_flush_pipe_pad;
  wire [11:0] wb_reg_replay_shl;
  wire [19:0] wb_reg_replay_pad;
  wire [8:0] id_reg_pause_shl;
  wire [19:0] id_reg_pause_pad;
  wire [3:0] wb_ctrl_rxs1_shl;
  wire [19:0] wb_ctrl_rxs1_pad;
  wire [17:0] ex_ctrl_rxs2_shl;
  wire [19:0] ex_ctrl_rxs2_pad;
  wire [1:0] ex_reg_replay_shl;
  wire [19:0] ex_reg_replay_pad;
  wire [7:0] mem_ctrl_div_shl;
  wire [19:0] mem_ctrl_div_pad;
  wire [12:0] wb_ctrl_wfd_shl;
  wire [19:0] wb_ctrl_wfd_pad;
  wire [12:0] wb_ctrl_mem_shl;
  wire [19:0] wb_ctrl_mem_pad;
  wire [19:0] wb_reg_flush_pipe_shl;
  wire [19:0] wb_reg_flush_pipe_pad;
  wire [8:0] mem_reg_rvc_shl;
  wire [19:0] mem_reg_rvc_pad;
  wire [8:0] mem_reg_xcpt_interrupt_shl;
  wire [19:0] mem_reg_xcpt_interrupt_pad;
  wire [3:0] ex_ctrl_mem_shl;
  wire [19:0] ex_ctrl_mem_pad;
  wire [10:0] ex_ctrl_sel_alu2_shl;
  wire [19:0] ex_ctrl_sel_alu2_pad;
  wire [4:0] id_reg_fence_shl;
  wire [19:0] id_reg_fence_pad;
  wire [14:0] mem_ctrl_wxd_shl;
  wire [19:0] mem_ctrl_wxd_pad;
  wire [2:0] mem_reg_xcpt_shl;
  wire [19:0] mem_reg_xcpt_pad;
  wire [19:0] ex_reg_valid_shl;
  wire [19:0] ex_reg_valid_pad;
  wire [14:0] ex_ctrl_div_shl;
  wire [19:0] ex_ctrl_div_pad;
  wire [5:0] ex_ctrl_wfd_shl;
  wire [19:0] ex_ctrl_wfd_pad;
  wire [4:0] wb_ctrl_rfs1_shl;
  wire [19:0] wb_ctrl_rfs1_pad;
  wire [7:0] mem_ctrl_fp_shl;
  wire [19:0] mem_ctrl_fp_pad;
  wire [11:0] mem_reg_sfence_shl;
  wire [19:0] mem_reg_sfence_pad;
  wire [12:0] wb_ctrl_div_shl;
  wire [19:0] wb_ctrl_div_pad;
  wire [9:0] mem_reg_replay_shl;
  wire [19:0] mem_reg_replay_pad;
  wire [14:0] ex_reg_rvc_shl;
  wire [19:0] ex_reg_rvc_pad;
  wire [6:0] blocked_shl;
  wire [19:0] blocked_pad;
  wire [5:0] mem_reg_valid_shl;
  wire [19:0] mem_reg_valid_pad;
  wire [16:0] mem_ctrl_jalr_shl;
  wire [19:0] mem_ctrl_jalr_pad;
  wire [8:0] wb_ctrl_wxd_shl;
  wire [19:0] wb_ctrl_wxd_pad;
  wire [17:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [17:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [9:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [10:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [15:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire  mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [10:0] ex_reg_rs_lsb_0_shl;
  wire [19:0] ex_reg_rs_lsb_0_pad;
  wire [10:0] ex_reg_rs_lsb_1_shl;
  wire [19:0] ex_reg_rs_lsb_1_pad;
  wire [13:0] ex_reg_rs_bypass_0_shl;
  wire [19:0] ex_reg_rs_bypass_0_pad;
  wire [13:0] ex_reg_rs_bypass_1_shl;
  wire [19:0] ex_reg_rs_bypass_1_pad;
  wire [19:0] Rocket_xor32;
  wire [19:0] Rocket_xor15;
  wire [19:0] Rocket_xor33;
  wire [19:0] Rocket_xor34;
  wire [19:0] Rocket_xor16;
  wire [19:0] Rocket_xor7;
  wire [19:0] Rocket_xor36;
  wire [19:0] Rocket_xor17;
  wire [19:0] Rocket_xor37;
  wire [19:0] Rocket_xor38;
  wire [19:0] Rocket_xor18;
  wire [19:0] Rocket_xor8;
  wire [19:0] Rocket_xor3;
  wire [19:0] Rocket_xor40;
  wire [19:0] Rocket_xor19;
  wire [19:0] Rocket_xor41;
  wire [19:0] Rocket_xor42;
  wire [19:0] Rocket_xor20;
  wire [19:0] Rocket_xor9;
  wire [19:0] Rocket_xor43;
  wire [19:0] Rocket_xor44;
  wire [19:0] Rocket_xor21;
  wire [19:0] Rocket_xor45;
  wire [19:0] Rocket_xor46;
  wire [19:0] Rocket_xor22;
  wire [19:0] Rocket_xor10;
  wire [19:0] Rocket_xor4;
  wire [19:0] Rocket_xor1;
  wire [19:0] Rocket_xor48;
  wire [19:0] Rocket_xor23;
  wire [19:0] Rocket_xor49;
  wire [19:0] Rocket_xor50;
  wire [19:0] Rocket_xor24;
  wire [19:0] Rocket_xor11;
  wire [19:0] Rocket_xor51;
  wire [19:0] Rocket_xor52;
  wire [19:0] Rocket_xor25;
  wire [19:0] Rocket_xor53;
  wire [19:0] Rocket_xor54;
  wire [19:0] Rocket_xor26;
  wire [19:0] Rocket_xor12;
  wire [19:0] Rocket_xor5;
  wire [19:0] Rocket_xor56;
  wire [19:0] Rocket_xor27;
  wire [19:0] Rocket_xor57;
  wire [19:0] Rocket_xor58;
  wire [19:0] Rocket_xor28;
  wire [19:0] Rocket_xor13;
  wire [19:0] Rocket_xor59;
  wire [19:0] Rocket_xor60;
  wire [19:0] Rocket_xor29;
  wire [19:0] Rocket_xor61;
  wire [19:0] Rocket_xor62;
  wire [19:0] Rocket_xor30;
  wire [19:0] Rocket_xor14;
  wire [19:0] Rocket_xor6;
  wire [19:0] Rocket_xor2;
  wire [19:0] Rocket_xor0;
  wire [29:0] alu_sum;
  wire [29:0] csr_sum;
  wire [29:0] div_sum;
  wire [29:0] bpu_sum;
  wire [29:0] ibuf_sum;
  wire [29:0] PlusArgTimeout_sum;
  wire  alu_metaAssert_wire;
  wire  div_metaAssert_wire;
  wire  bpu_metaAssert_wire;
  wire  PlusArgTimeout_metaAssert_wire;
  wire  ibuf_metaAssert_wire;
  wire  csr_metaAssert_wire;
  wire  Rocket_or4;
  wire  Rocket_or1;
  wire  Rocket_or6;
  wire  Rocket_or2;
  wire  Rocket_or0;
  reg  Rocket_metaAssert;
  reg [31:0] _RAND_112;
  IBuf ibuf ( // @[RocketCore.scala 248:20]
    .clock(ibuf_clock),
    .reset(ibuf_reset),
    .io_imem_ready(ibuf_io_imem_ready),
    .io_imem_valid(ibuf_io_imem_valid),
    .io_imem_bits_btb_taken(ibuf_io_imem_bits_btb_taken),
    .io_imem_bits_btb_bridx(ibuf_io_imem_bits_btb_bridx),
    .io_imem_bits_btb_entry(ibuf_io_imem_bits_btb_entry),
    .io_imem_bits_btb_bht_history(ibuf_io_imem_bits_btb_bht_history),
    .io_imem_bits_pc(ibuf_io_imem_bits_pc),
    .io_imem_bits_data(ibuf_io_imem_bits_data),
    .io_imem_bits_xcpt_pf_inst(ibuf_io_imem_bits_xcpt_pf_inst),
    .io_imem_bits_xcpt_ae_inst(ibuf_io_imem_bits_xcpt_ae_inst),
    .io_imem_bits_replay(ibuf_io_imem_bits_replay),
    .io_kill(ibuf_io_kill),
    .io_pc(ibuf_io_pc),
    .io_btb_resp_entry(ibuf_io_btb_resp_entry),
    .io_btb_resp_bht_history(ibuf_io_btb_resp_bht_history),
    .io_inst_0_ready(ibuf_io_inst_0_ready),
    .io_inst_0_valid(ibuf_io_inst_0_valid),
    .io_inst_0_bits_xcpt0_pf_inst(ibuf_io_inst_0_bits_xcpt0_pf_inst),
    .io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),
    .io_inst_0_bits_xcpt1_pf_inst(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .io_inst_0_bits_xcpt1_ae_inst(ibuf_io_inst_0_bits_xcpt1_ae_inst),
    .io_inst_0_bits_replay(ibuf_io_inst_0_bits_replay),
    .io_inst_0_bits_rvc(ibuf_io_inst_0_bits_rvc),
    .io_inst_0_bits_inst_bits(ibuf_io_inst_0_bits_inst_bits),
    .io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
    .io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
    .io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
    .io_inst_0_bits_inst_rs3(ibuf_io_inst_0_bits_inst_rs3),
    .io_inst_0_bits_raw(ibuf_io_inst_0_bits_raw),
    .io_covSum(ibuf_io_covSum),
    .metaAssert(ibuf_metaAssert),
    .metaReset(ibuf_metaReset)
  );
  CSRFile csr ( // @[RocketCore.scala 276:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_ungated_clock(csr_io_ungated_clock),
    .io_interrupts_debug(csr_io_interrupts_debug),
    .io_interrupts_mtip(csr_io_interrupts_mtip),
    .io_interrupts_msip(csr_io_interrupts_msip),
    .io_interrupts_meip(csr_io_interrupts_meip),
    .io_interrupts_seip(csr_io_interrupts_seip),
    .io_hartid(csr_io_hartid),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_decode_0_csr(csr_io_decode_0_csr),
    .io_decode_0_fp_illegal(csr_io_decode_0_fp_illegal),
    .io_decode_0_fp_csr(csr_io_decode_0_fp_csr),
    .io_decode_0_read_illegal(csr_io_decode_0_read_illegal),
    .io_decode_0_write_illegal(csr_io_decode_0_write_illegal),
    .io_decode_0_write_flush(csr_io_decode_0_write_flush),
    .io_decode_0_system_illegal(csr_io_decode_0_system_illegal),
    .io_csr_stall(csr_io_csr_stall),
    .io_eret(csr_io_eret),
    .io_singleStep(csr_io_singleStep),
    .io_status_debug(csr_io_status_debug),
    .io_status_cease(csr_io_status_cease),
    .io_status_wfi(csr_io_status_wfi),
    .io_status_isa(csr_io_status_isa),
    .io_status_dprv(csr_io_status_dprv),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero2(csr_io_status_zero2),
    .io_status_sxl(csr_io_status_sxl),
    .io_status_uxl(csr_io_status_uxl),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_tsr(csr_io_status_tsr),
    .io_status_tw(csr_io_status_tw),
    .io_status_tvm(csr_io_status_tvm),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_sum(csr_io_status_sum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_vs(csr_io_status_vs),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_ptbr_mode(csr_io_ptbr_mode),
    .io_ptbr_ppn(csr_io_ptbr_ppn),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_cause(csr_io_cause),
    .io_pc(csr_io_pc),
    .io_tval(csr_io_tval),
    .io_time(csr_io_time),
    .io_fcsr_rm(csr_io_fcsr_rm),
    .io_fcsr_flags_valid(csr_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(csr_io_fcsr_flags_bits),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_bp_0_control_action(csr_io_bp_0_control_action),
    .io_bp_0_control_tmatch(csr_io_bp_0_control_tmatch),
    .io_bp_0_control_m(csr_io_bp_0_control_m),
    .io_bp_0_control_s(csr_io_bp_0_control_s),
    .io_bp_0_control_u(csr_io_bp_0_control_u),
    .io_bp_0_control_x(csr_io_bp_0_control_x),
    .io_bp_0_control_w(csr_io_bp_0_control_w),
    .io_bp_0_control_r(csr_io_bp_0_control_r),
    .io_bp_0_address(csr_io_bp_0_address),
    .io_pmp_0_cfg_l(csr_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(csr_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(csr_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(csr_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(csr_io_pmp_0_cfg_r),
    .io_pmp_0_addr(csr_io_pmp_0_addr),
    .io_pmp_0_mask(csr_io_pmp_0_mask),
    .io_pmp_1_cfg_l(csr_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(csr_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(csr_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(csr_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(csr_io_pmp_1_cfg_r),
    .io_pmp_1_addr(csr_io_pmp_1_addr),
    .io_pmp_1_mask(csr_io_pmp_1_mask),
    .io_pmp_2_cfg_l(csr_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(csr_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(csr_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(csr_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(csr_io_pmp_2_cfg_r),
    .io_pmp_2_addr(csr_io_pmp_2_addr),
    .io_pmp_2_mask(csr_io_pmp_2_mask),
    .io_pmp_3_cfg_l(csr_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(csr_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(csr_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(csr_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(csr_io_pmp_3_cfg_r),
    .io_pmp_3_addr(csr_io_pmp_3_addr),
    .io_pmp_3_mask(csr_io_pmp_3_mask),
    .io_pmp_4_cfg_l(csr_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(csr_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(csr_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(csr_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(csr_io_pmp_4_cfg_r),
    .io_pmp_4_addr(csr_io_pmp_4_addr),
    .io_pmp_4_mask(csr_io_pmp_4_mask),
    .io_pmp_5_cfg_l(csr_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(csr_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(csr_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(csr_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(csr_io_pmp_5_cfg_r),
    .io_pmp_5_addr(csr_io_pmp_5_addr),
    .io_pmp_5_mask(csr_io_pmp_5_mask),
    .io_pmp_6_cfg_l(csr_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(csr_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(csr_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(csr_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(csr_io_pmp_6_cfg_r),
    .io_pmp_6_addr(csr_io_pmp_6_addr),
    .io_pmp_6_mask(csr_io_pmp_6_mask),
    .io_pmp_7_cfg_l(csr_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(csr_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(csr_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(csr_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(csr_io_pmp_7_cfg_r),
    .io_pmp_7_addr(csr_io_pmp_7_addr),
    .io_pmp_7_mask(csr_io_pmp_7_mask),
    .io_inst_0(csr_io_inst_0),
    .io_trace_0_valid(csr_io_trace_0_valid),
    .io_trace_0_iaddr(csr_io_trace_0_iaddr),
    .io_trace_0_insn(csr_io_trace_0_insn),
    .io_trace_0_exception(csr_io_trace_0_exception),
    .io_customCSRs_0_value(csr_io_customCSRs_0_value),
    .io_covSum(csr_io_covSum),
    .metaAssert(csr_metaAssert),
    .metaReset(csr_metaReset)
  );
  BreakpointUnit bpu ( // @[RocketCore.scala 317:19]
    .io_status_debug(bpu_io_status_debug),
    .io_status_prv(bpu_io_status_prv),
    .io_bp_0_control_action(bpu_io_bp_0_control_action),
    .io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),
    .io_bp_0_control_m(bpu_io_bp_0_control_m),
    .io_bp_0_control_s(bpu_io_bp_0_control_s),
    .io_bp_0_control_u(bpu_io_bp_0_control_u),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_pc(bpu_io_pc),
    .io_ea(bpu_io_ea),
    .io_xcpt_if(bpu_io_xcpt_if),
    .io_xcpt_ld(bpu_io_xcpt_ld),
    .io_xcpt_st(bpu_io_xcpt_st),
    .io_debug_if(bpu_io_debug_if),
    .io_debug_ld(bpu_io_debug_ld),
    .io_debug_st(bpu_io_debug_st),
    .io_covSum(bpu_io_covSum),
    .metaAssert(bpu_metaAssert)
  );
  ALU alu ( // @[RocketCore.scala 377:19]
    .io_dw(alu_io_dw),
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out),
    .io_covSum(alu_io_covSum),
    .metaAssert(alu_metaAssert)
  );
  MulDiv div ( // @[RocketCore.scala 401:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_req_bits_fn(div_io_req_bits_fn),
    .io_req_bits_dw(div_io_req_bits_dw),
    .io_req_bits_in1(div_io_req_bits_in1),
    .io_req_bits_in2(div_io_req_bits_in2),
    .io_req_bits_tag(div_io_req_bits_tag),
    .io_kill(div_io_kill),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag),
    .io_covSum(div_io_covSum),
    .metaAssert(div_metaAssert),
    .metaReset(div_metaReset)
  );
  PlusArgTimeout PlusArgTimeout ( // @[PlusArg.scala 89:11]
    .io_covSum(PlusArgTimeout_io_covSum),
    .metaAssert(PlusArgTimeout_metaAssert)
  );
  assign _T_815__T_820_addr = ~id_raddr1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_815__T_820_data = _T_815[_T_815__T_820_addr]; // @[RocketCore.scala 1014:15]
  `else
  assign _T_815__T_820_data = _T_815__T_820_addr >= 5'h1f ? _RAND_1[63:0] : _T_815[_T_815__T_820_addr]; // @[RocketCore.scala 1014:15]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_815__T_826_addr = ~id_raddr2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_815__T_826_data = _T_815[_T_815__T_826_addr]; // @[RocketCore.scala 1014:15]
  `else
  assign _T_815__T_826_data = _T_815__T_826_addr >= 5'h1f ? _RAND_2[63:0] : _T_815[_T_815__T_826_addr]; // @[RocketCore.scala 1014:15]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_815__T_1524_data = _T_1515 ? io_dmem_resp_bits_data : _T_1520;
  assign _T_815__T_1524_addr = ~rf_waddr;
  assign _T_815__T_1524_mask = 1'h1;
  assign _T_815__T_1524_en = rf_wen & _T_1521;
  assign replay_wb_common = io_dmem_s2_nack | wb_reg_replay; // @[RocketCore.scala 629:42]
  assign _T_1465 = wb_reg_valid & wb_ctrl_mem; // @[RocketCore.scala 607:19]
  assign _T_1466 = _T_1465 & io_dmem_s2_xcpt_ma_st; // @[RocketCore.scala 607:34]
  assign _T_1477 = wb_reg_xcpt | _T_1466; // @[RocketCore.scala 974:26]
  assign _T_1468 = _T_1465 & io_dmem_s2_xcpt_ma_ld; // @[RocketCore.scala 608:34]
  assign _T_1478 = _T_1477 | _T_1468; // @[RocketCore.scala 974:26]
  assign _T_1470 = _T_1465 & io_dmem_s2_xcpt_pf_st; // @[RocketCore.scala 609:34]
  assign _T_1479 = _T_1478 | _T_1470; // @[RocketCore.scala 974:26]
  assign _T_1472 = _T_1465 & io_dmem_s2_xcpt_pf_ld; // @[RocketCore.scala 610:34]
  assign _T_1480 = _T_1479 | _T_1472; // @[RocketCore.scala 974:26]
  assign _T_1474 = _T_1465 & io_dmem_s2_xcpt_ae_st; // @[RocketCore.scala 611:34]
  assign _T_1481 = _T_1480 | _T_1474; // @[RocketCore.scala 974:26]
  assign _T_1476 = _T_1465 & io_dmem_s2_xcpt_ae_ld; // @[RocketCore.scala 612:34]
  assign wb_xcpt = _T_1481 | _T_1476; // @[RocketCore.scala 974:26]
  assign _T_1503 = replay_wb_common | wb_xcpt; // @[RocketCore.scala 632:27]
  assign _T_1504 = _T_1503 | csr_io_eret; // @[RocketCore.scala 632:38]
  assign take_pc_wb = _T_1504 | wb_reg_flush_pipe; // @[RocketCore.scala 632:53]
  assign _T_1149 = ex_reg_valid | ex_reg_replay; // @[RocketCore.scala 482:34]
  assign ex_pc_valid = _T_1149 | ex_reg_xcpt_interrupt; // @[RocketCore.scala 482:51]
  assign _T_1305 = mem_ctrl_jalr | mem_reg_sfence; // @[RocketCore.scala 505:36]
  assign a = mem_reg_wdata[63:39]; // @[RocketCore.scala 988:23]
  assign _T_1307 = $signed(a) == 25'sh0; // @[RocketCore.scala 989:21]
  assign _T_1308 = $signed(a) == -25'sh1; // @[RocketCore.scala 989:34]
  assign _T_1309 = _T_1307 | _T_1308; // @[RocketCore.scala 989:29]
  assign msb = _T_1309 ? mem_reg_wdata[39] : ~mem_reg_wdata[38]; // @[RocketCore.scala 989:18]
  assign _T_1315 = {msb,mem_reg_wdata[38:0]}; // @[RocketCore.scala 505:106]
  assign _T_1175 = mem_ctrl_branch & mem_br_taken; // @[RocketCore.scala 502:25]
  assign _T_1178 = mem_reg_inst[31]; // @[RocketCore.scala 1036:53]
  assign _T_1233 = mem_reg_inst[31]; // @[Cat.scala 29:58]
  assign _T_1232 = {11{_T_1178}}; // @[Cat.scala 29:58]
  assign _T_1230 = {8{_T_1178}}; // @[Cat.scala 29:58]
  assign _T_1229 = mem_reg_inst[7]; // @[Cat.scala 29:58]
  assign _T_1237 = {_T_1233,_T_1232,_T_1230,_T_1229,mem_reg_inst[30:25],mem_reg_inst[11:8],1'h0}; // @[RocketCore.scala 1050:53]
  assign _T_1292 = mem_reg_inst[19:12]; // @[Cat.scala 29:58]
  assign _T_1291 = mem_reg_inst[20]; // @[Cat.scala 29:58]
  assign _T_1299 = {_T_1233,_T_1232,_T_1292,_T_1291,mem_reg_inst[30:25],mem_reg_inst[24:21],1'h0}; // @[RocketCore.scala 1050:53]
  assign _T_1300 = mem_reg_rvc ? $signed(4'sh2) : $signed(4'sh4); // @[RocketCore.scala 504:8]
  assign _T_1301 = mem_ctrl_jal ? $signed(_T_1299) : $signed({{28{_T_1300[3]}},_T_1300}); // @[RocketCore.scala 503:8]
  assign _T_1302 = _T_1175 ? $signed(_T_1237) : $signed(_T_1301); // @[RocketCore.scala 502:8]
  assign _GEN_248 = {{8{_T_1302[31]}},_T_1302}; // @[RocketCore.scala 501:41]
  assign mem_br_target = $signed(mem_reg_pc) + $signed(_GEN_248); // @[RocketCore.scala 501:41]
  assign _T_1316 = _T_1305 ? $signed(_T_1315) : $signed(mem_br_target); // @[RocketCore.scala 505:21]
  assign mem_npc = $signed(_T_1316) & -40'sh2; // @[RocketCore.scala 505:141]
  assign _T_1319 = mem_npc != ex_reg_pc; // @[RocketCore.scala 507:30]
  assign _T_1320 = ibuf_io_inst_0_valid | ibuf_io_imem_valid; // @[RocketCore.scala 508:31]
  assign _T_1321 = mem_npc != ibuf_io_pc; // @[RocketCore.scala 508:62]
  assign _T_1322 = _T_1320 ? _T_1321 : 1'h1; // @[RocketCore.scala 508:8]
  assign mem_wrong_npc = ex_pc_valid ? _T_1319 : _T_1322; // @[RocketCore.scala 507:8]
  assign _T_1338 = mem_wrong_npc | mem_reg_sfence; // @[RocketCore.scala 515:54]
  assign take_pc_mem = mem_reg_valid & _T_1338; // @[RocketCore.scala 515:32]
  assign take_pc_mem_wb = take_pc_wb | take_pc_mem; // @[RocketCore.scala 244:35]
  assign _T_3 = ibuf_io_inst_0_bits_inst_bits & 32'hfe00707f; // @[Decode.scala 14:65]
  assign _T_4 = _T_3 == 32'h2000033; // @[Decode.scala 14:121]
  assign _T_6 = _T_3 == 32'h2001033; // @[Decode.scala 14:121]
  assign _T_8 = _T_3 == 32'h2003033; // @[Decode.scala 14:121]
  assign _T_10 = _T_3 == 32'h2002033; // @[Decode.scala 14:121]
  assign _T_12 = _T_3 == 32'h2004033; // @[Decode.scala 14:121]
  assign _T_14 = _T_3 == 32'h2005033; // @[Decode.scala 14:121]
  assign _T_16 = _T_3 == 32'h2006033; // @[Decode.scala 14:121]
  assign _T_18 = _T_3 == 32'h2007033; // @[Decode.scala 14:121]
  assign _T_20 = _T_3 == 32'h200003b; // @[Decode.scala 14:121]
  assign _T_22 = _T_3 == 32'h200403b; // @[Decode.scala 14:121]
  assign _T_24 = _T_3 == 32'h200503b; // @[Decode.scala 14:121]
  assign _T_26 = _T_3 == 32'h200603b; // @[Decode.scala 14:121]
  assign _T_28 = _T_3 == 32'h200703b; // @[Decode.scala 14:121]
  assign _T_29 = ibuf_io_inst_0_bits_inst_bits & 32'hf800707f; // @[Decode.scala 14:65]
  assign _T_30 = _T_29 == 32'h202f; // @[Decode.scala 14:121]
  assign _T_32 = _T_29 == 32'h2000202f; // @[Decode.scala 14:121]
  assign _T_34 = _T_29 == 32'h800202f; // @[Decode.scala 14:121]
  assign _T_36 = _T_29 == 32'h6000202f; // @[Decode.scala 14:121]
  assign _T_38 = _T_29 == 32'h4000202f; // @[Decode.scala 14:121]
  assign _T_40 = _T_29 == 32'h8000202f; // @[Decode.scala 14:121]
  assign _T_42 = _T_29 == 32'hc000202f; // @[Decode.scala 14:121]
  assign _T_44 = _T_29 == 32'ha000202f; // @[Decode.scala 14:121]
  assign _T_46 = _T_29 == 32'he000202f; // @[Decode.scala 14:121]
  assign _T_47 = ibuf_io_inst_0_bits_inst_bits & 32'hf9f0707f; // @[Decode.scala 14:65]
  assign _T_48 = _T_47 == 32'h1000202f; // @[Decode.scala 14:121]
  assign _T_50 = _T_29 == 32'h1800202f; // @[Decode.scala 14:121]
  assign _T_52 = _T_29 == 32'h302f; // @[Decode.scala 14:121]
  assign _T_54 = _T_29 == 32'h800302f; // @[Decode.scala 14:121]
  assign _T_56 = _T_29 == 32'h2000302f; // @[Decode.scala 14:121]
  assign _T_58 = _T_29 == 32'h6000302f; // @[Decode.scala 14:121]
  assign _T_60 = _T_29 == 32'h4000302f; // @[Decode.scala 14:121]
  assign _T_62 = _T_29 == 32'h8000302f; // @[Decode.scala 14:121]
  assign _T_64 = _T_29 == 32'hc000302f; // @[Decode.scala 14:121]
  assign _T_66 = _T_29 == 32'ha000302f; // @[Decode.scala 14:121]
  assign _T_68 = _T_29 == 32'he000302f; // @[Decode.scala 14:121]
  assign _T_70 = _T_47 == 32'h1000302f; // @[Decode.scala 14:121]
  assign _T_72 = _T_29 == 32'h1800302f; // @[Decode.scala 14:121]
  assign _T_74 = _T_3 == 32'h20000053; // @[Decode.scala 14:121]
  assign _T_76 = _T_3 == 32'h20002053; // @[Decode.scala 14:121]
  assign _T_78 = _T_3 == 32'h20001053; // @[Decode.scala 14:121]
  assign _T_80 = _T_3 == 32'h28000053; // @[Decode.scala 14:121]
  assign _T_82 = _T_3 == 32'h28001053; // @[Decode.scala 14:121]
  assign _T_83 = ibuf_io_inst_0_bits_inst_bits & 32'hfe00007f; // @[Decode.scala 14:65]
  assign _T_84 = _T_83 == 32'h53; // @[Decode.scala 14:121]
  assign _T_86 = _T_83 == 32'h8000053; // @[Decode.scala 14:121]
  assign _T_88 = _T_83 == 32'h10000053; // @[Decode.scala 14:121]
  assign _T_89 = ibuf_io_inst_0_bits_inst_bits & 32'h600007f; // @[Decode.scala 14:65]
  assign _T_90 = _T_89 == 32'h43; // @[Decode.scala 14:121]
  assign _T_92 = _T_89 == 32'h47; // @[Decode.scala 14:121]
  assign _T_94 = _T_89 == 32'h4f; // @[Decode.scala 14:121]
  assign _T_96 = _T_89 == 32'h4b; // @[Decode.scala 14:121]
  assign _T_97 = ibuf_io_inst_0_bits_inst_bits & 32'hfff0707f; // @[Decode.scala 14:65]
  assign _T_98 = _T_97 == 32'he0001053; // @[Decode.scala 14:121]
  assign _T_100 = _T_97 == 32'he0000053; // @[Decode.scala 14:121]
  assign _T_101 = ibuf_io_inst_0_bits_inst_bits & 32'hfff0007f; // @[Decode.scala 14:65]
  assign _T_102 = _T_101 == 32'hc0000053; // @[Decode.scala 14:121]
  assign _T_104 = _T_101 == 32'hc0100053; // @[Decode.scala 14:121]
  assign _T_106 = _T_3 == 32'ha0002053; // @[Decode.scala 14:121]
  assign _T_108 = _T_3 == 32'ha0001053; // @[Decode.scala 14:121]
  assign _T_110 = _T_3 == 32'ha0000053; // @[Decode.scala 14:121]
  assign _T_112 = _T_97 == 32'hf0000053; // @[Decode.scala 14:121]
  assign _T_114 = _T_101 == 32'hd0000053; // @[Decode.scala 14:121]
  assign _T_116 = _T_101 == 32'hd0100053; // @[Decode.scala 14:121]
  assign _T_117 = ibuf_io_inst_0_bits_inst_bits & 32'h707f; // @[Decode.scala 14:65]
  assign _T_118 = _T_117 == 32'h2007; // @[Decode.scala 14:121]
  assign _T_120 = _T_117 == 32'h2027; // @[Decode.scala 14:121]
  assign _T_122 = _T_83 == 32'h18000053; // @[Decode.scala 14:121]
  assign _T_124 = _T_101 == 32'h58000053; // @[Decode.scala 14:121]
  assign _T_126 = _T_101 == 32'hc0200053; // @[Decode.scala 14:121]
  assign _T_128 = _T_101 == 32'hc0300053; // @[Decode.scala 14:121]
  assign _T_130 = _T_101 == 32'hd0200053; // @[Decode.scala 14:121]
  assign _T_132 = _T_101 == 32'hd0300053; // @[Decode.scala 14:121]
  assign _T_134 = _T_101 == 32'h40100053; // @[Decode.scala 14:121]
  assign _T_136 = _T_101 == 32'h42000053; // @[Decode.scala 14:121]
  assign _T_138 = _T_3 == 32'h22000053; // @[Decode.scala 14:121]
  assign _T_140 = _T_3 == 32'h22002053; // @[Decode.scala 14:121]
  assign _T_142 = _T_3 == 32'h22001053; // @[Decode.scala 14:121]
  assign _T_144 = _T_3 == 32'h2a000053; // @[Decode.scala 14:121]
  assign _T_146 = _T_3 == 32'h2a001053; // @[Decode.scala 14:121]
  assign _T_148 = _T_83 == 32'h2000053; // @[Decode.scala 14:121]
  assign _T_150 = _T_83 == 32'ha000053; // @[Decode.scala 14:121]
  assign _T_152 = _T_83 == 32'h12000053; // @[Decode.scala 14:121]
  assign _T_154 = _T_89 == 32'h2000043; // @[Decode.scala 14:121]
  assign _T_156 = _T_89 == 32'h2000047; // @[Decode.scala 14:121]
  assign _T_158 = _T_89 == 32'h200004f; // @[Decode.scala 14:121]
  assign _T_160 = _T_89 == 32'h200004b; // @[Decode.scala 14:121]
  assign _T_162 = _T_97 == 32'he2001053; // @[Decode.scala 14:121]
  assign _T_164 = _T_101 == 32'hc2000053; // @[Decode.scala 14:121]
  assign _T_166 = _T_101 == 32'hc2100053; // @[Decode.scala 14:121]
  assign _T_168 = _T_3 == 32'ha2002053; // @[Decode.scala 14:121]
  assign _T_170 = _T_3 == 32'ha2001053; // @[Decode.scala 14:121]
  assign _T_172 = _T_3 == 32'ha2000053; // @[Decode.scala 14:121]
  assign _T_174 = _T_101 == 32'hd2000053; // @[Decode.scala 14:121]
  assign _T_176 = _T_101 == 32'hd2100053; // @[Decode.scala 14:121]
  assign _T_178 = _T_117 == 32'h3007; // @[Decode.scala 14:121]
  assign _T_180 = _T_117 == 32'h3027; // @[Decode.scala 14:121]
  assign _T_182 = _T_83 == 32'h1a000053; // @[Decode.scala 14:121]
  assign _T_184 = _T_101 == 32'h5a000053; // @[Decode.scala 14:121]
  assign _T_186 = _T_97 == 32'he2000053; // @[Decode.scala 14:121]
  assign _T_188 = _T_101 == 32'hc2200053; // @[Decode.scala 14:121]
  assign _T_190 = _T_101 == 32'hc2300053; // @[Decode.scala 14:121]
  assign _T_192 = _T_97 == 32'hf2000053; // @[Decode.scala 14:121]
  assign _T_194 = _T_101 == 32'hd2200053; // @[Decode.scala 14:121]
  assign _T_196 = _T_101 == 32'hd2300053; // @[Decode.scala 14:121]
  assign _T_198 = _T_117 == 32'h3003; // @[Decode.scala 14:121]
  assign _T_200 = _T_117 == 32'h6003; // @[Decode.scala 14:121]
  assign _T_202 = _T_117 == 32'h3023; // @[Decode.scala 14:121]
  assign _T_203 = ibuf_io_inst_0_bits_inst_bits & 32'hfc00707f; // @[Decode.scala 14:65]
  assign _T_204 = _T_203 == 32'h1013; // @[Decode.scala 14:121]
  assign _T_206 = _T_203 == 32'h5013; // @[Decode.scala 14:121]
  assign _T_208 = _T_203 == 32'h40005013; // @[Decode.scala 14:121]
  assign _T_210 = _T_117 == 32'h1b; // @[Decode.scala 14:121]
  assign _T_212 = _T_3 == 32'h101b; // @[Decode.scala 14:121]
  assign _T_214 = _T_3 == 32'h501b; // @[Decode.scala 14:121]
  assign _T_216 = _T_3 == 32'h4000501b; // @[Decode.scala 14:121]
  assign _T_218 = _T_3 == 32'h3b; // @[Decode.scala 14:121]
  assign _T_220 = _T_3 == 32'h4000003b; // @[Decode.scala 14:121]
  assign _T_222 = _T_3 == 32'h103b; // @[Decode.scala 14:121]
  assign _T_224 = _T_3 == 32'h503b; // @[Decode.scala 14:121]
  assign _T_226 = _T_3 == 32'h4000503b; // @[Decode.scala 14:121]
  assign _T_227 = ibuf_io_inst_0_bits_inst_bits & 32'hfe007fff; // @[Decode.scala 14:65]
  assign _T_228 = _T_227 == 32'h12000073; // @[Decode.scala 14:121]
  assign _T_229 = ibuf_io_inst_0_bits_inst_bits == 32'h10200073; // @[Decode.scala 14:121]
  assign _T_230 = ibuf_io_inst_0_bits_inst_bits == 32'h7b200073; // @[Decode.scala 14:121]
  assign _T_232 = _T_117 == 32'h100f; // @[Decode.scala 14:121]
  assign _T_234 = _T_117 == 32'h1063; // @[Decode.scala 14:121]
  assign _T_236 = _T_117 == 32'h63; // @[Decode.scala 14:121]
  assign _T_238 = _T_117 == 32'h4063; // @[Decode.scala 14:121]
  assign _T_240 = _T_117 == 32'h6063; // @[Decode.scala 14:121]
  assign _T_242 = _T_117 == 32'h5063; // @[Decode.scala 14:121]
  assign _T_244 = _T_117 == 32'h7063; // @[Decode.scala 14:121]
  assign _T_245 = ibuf_io_inst_0_bits_inst_bits & 32'h7f; // @[Decode.scala 14:65]
  assign _T_246 = _T_245 == 32'h6f; // @[Decode.scala 14:121]
  assign _T_248 = _T_117 == 32'h67; // @[Decode.scala 14:121]
  assign _T_250 = _T_245 == 32'h17; // @[Decode.scala 14:121]
  assign _T_252 = _T_117 == 32'h3; // @[Decode.scala 14:121]
  assign _T_254 = _T_117 == 32'h1003; // @[Decode.scala 14:121]
  assign _T_256 = _T_117 == 32'h2003; // @[Decode.scala 14:121]
  assign _T_258 = _T_117 == 32'h4003; // @[Decode.scala 14:121]
  assign _T_260 = _T_117 == 32'h5003; // @[Decode.scala 14:121]
  assign _T_262 = _T_117 == 32'h23; // @[Decode.scala 14:121]
  assign _T_264 = _T_117 == 32'h1023; // @[Decode.scala 14:121]
  assign _T_266 = _T_117 == 32'h2023; // @[Decode.scala 14:121]
  assign _T_268 = _T_245 == 32'h37; // @[Decode.scala 14:121]
  assign _T_270 = _T_117 == 32'h13; // @[Decode.scala 14:121]
  assign _T_272 = _T_117 == 32'h2013; // @[Decode.scala 14:121]
  assign _T_274 = _T_117 == 32'h3013; // @[Decode.scala 14:121]
  assign _T_276 = _T_117 == 32'h7013; // @[Decode.scala 14:121]
  assign _T_278 = _T_117 == 32'h6013; // @[Decode.scala 14:121]
  assign _T_280 = _T_117 == 32'h4013; // @[Decode.scala 14:121]
  assign _T_282 = _T_3 == 32'h33; // @[Decode.scala 14:121]
  assign _T_284 = _T_3 == 32'h40000033; // @[Decode.scala 14:121]
  assign _T_286 = _T_3 == 32'h2033; // @[Decode.scala 14:121]
  assign _T_288 = _T_3 == 32'h3033; // @[Decode.scala 14:121]
  assign _T_290 = _T_3 == 32'h7033; // @[Decode.scala 14:121]
  assign _T_292 = _T_3 == 32'h6033; // @[Decode.scala 14:121]
  assign _T_294 = _T_3 == 32'h4033; // @[Decode.scala 14:121]
  assign _T_296 = _T_3 == 32'h1033; // @[Decode.scala 14:121]
  assign _T_298 = _T_3 == 32'h5033; // @[Decode.scala 14:121]
  assign _T_300 = _T_3 == 32'h40005033; // @[Decode.scala 14:121]
  assign _T_302 = _T_117 == 32'hf; // @[Decode.scala 14:121]
  assign _T_303 = ibuf_io_inst_0_bits_inst_bits == 32'h73; // @[Decode.scala 14:121]
  assign _T_304 = ibuf_io_inst_0_bits_inst_bits == 32'h100073; // @[Decode.scala 14:121]
  assign _T_305 = ibuf_io_inst_0_bits_inst_bits == 32'h30200073; // @[Decode.scala 14:121]
  assign _T_306 = ibuf_io_inst_0_bits_inst_bits == 32'h10500073; // @[Decode.scala 14:121]
  assign _T_307 = ibuf_io_inst_0_bits_inst_bits == 32'h30500073; // @[Decode.scala 14:121]
  assign _T_309 = _T_117 == 32'h1073; // @[Decode.scala 14:121]
  assign _T_311 = _T_117 == 32'h2073; // @[Decode.scala 14:121]
  assign _T_313 = _T_117 == 32'h3073; // @[Decode.scala 14:121]
  assign _T_315 = _T_117 == 32'h5073; // @[Decode.scala 14:121]
  assign _T_317 = _T_117 == 32'h6073; // @[Decode.scala 14:121]
  assign _T_319 = _T_117 == 32'h7073; // @[Decode.scala 14:121]
  assign _T_321 = _T_4 | _T_6; // @[Decode.scala 15:30]
  assign _T_322 = _T_321 | _T_8; // @[Decode.scala 15:30]
  assign _T_323 = _T_322 | _T_10; // @[Decode.scala 15:30]
  assign _T_324 = _T_323 | _T_12; // @[Decode.scala 15:30]
  assign _T_325 = _T_324 | _T_14; // @[Decode.scala 15:30]
  assign _T_326 = _T_325 | _T_16; // @[Decode.scala 15:30]
  assign _T_327 = _T_326 | _T_18; // @[Decode.scala 15:30]
  assign _T_328 = _T_327 | _T_20; // @[Decode.scala 15:30]
  assign _T_329 = _T_328 | _T_22; // @[Decode.scala 15:30]
  assign _T_330 = _T_329 | _T_24; // @[Decode.scala 15:30]
  assign _T_331 = _T_330 | _T_26; // @[Decode.scala 15:30]
  assign _T_332 = _T_331 | _T_28; // @[Decode.scala 15:30]
  assign _T_333 = _T_332 | _T_30; // @[Decode.scala 15:30]
  assign _T_334 = _T_333 | _T_32; // @[Decode.scala 15:30]
  assign _T_335 = _T_334 | _T_34; // @[Decode.scala 15:30]
  assign _T_336 = _T_335 | _T_36; // @[Decode.scala 15:30]
  assign _T_337 = _T_336 | _T_38; // @[Decode.scala 15:30]
  assign _T_338 = _T_337 | _T_40; // @[Decode.scala 15:30]
  assign _T_339 = _T_338 | _T_42; // @[Decode.scala 15:30]
  assign _T_340 = _T_339 | _T_44; // @[Decode.scala 15:30]
  assign _T_341 = _T_340 | _T_46; // @[Decode.scala 15:30]
  assign _T_342 = _T_341 | _T_48; // @[Decode.scala 15:30]
  assign _T_343 = _T_342 | _T_50; // @[Decode.scala 15:30]
  assign _T_344 = _T_343 | _T_52; // @[Decode.scala 15:30]
  assign _T_345 = _T_344 | _T_54; // @[Decode.scala 15:30]
  assign _T_346 = _T_345 | _T_56; // @[Decode.scala 15:30]
  assign _T_347 = _T_346 | _T_58; // @[Decode.scala 15:30]
  assign _T_348 = _T_347 | _T_60; // @[Decode.scala 15:30]
  assign _T_349 = _T_348 | _T_62; // @[Decode.scala 15:30]
  assign _T_350 = _T_349 | _T_64; // @[Decode.scala 15:30]
  assign _T_351 = _T_350 | _T_66; // @[Decode.scala 15:30]
  assign _T_352 = _T_351 | _T_68; // @[Decode.scala 15:30]
  assign _T_353 = _T_352 | _T_70; // @[Decode.scala 15:30]
  assign _T_354 = _T_353 | _T_72; // @[Decode.scala 15:30]
  assign _T_355 = _T_354 | _T_74; // @[Decode.scala 15:30]
  assign _T_356 = _T_355 | _T_76; // @[Decode.scala 15:30]
  assign _T_357 = _T_356 | _T_78; // @[Decode.scala 15:30]
  assign _T_358 = _T_357 | _T_80; // @[Decode.scala 15:30]
  assign _T_359 = _T_358 | _T_82; // @[Decode.scala 15:30]
  assign _T_360 = _T_359 | _T_84; // @[Decode.scala 15:30]
  assign _T_361 = _T_360 | _T_86; // @[Decode.scala 15:30]
  assign _T_362 = _T_361 | _T_88; // @[Decode.scala 15:30]
  assign _T_363 = _T_362 | _T_90; // @[Decode.scala 15:30]
  assign _T_364 = _T_363 | _T_92; // @[Decode.scala 15:30]
  assign _T_365 = _T_364 | _T_94; // @[Decode.scala 15:30]
  assign _T_366 = _T_365 | _T_96; // @[Decode.scala 15:30]
  assign _T_367 = _T_366 | _T_98; // @[Decode.scala 15:30]
  assign _T_368 = _T_367 | _T_100; // @[Decode.scala 15:30]
  assign _T_369 = _T_368 | _T_102; // @[Decode.scala 15:30]
  assign _T_370 = _T_369 | _T_104; // @[Decode.scala 15:30]
  assign _T_371 = _T_370 | _T_106; // @[Decode.scala 15:30]
  assign _T_372 = _T_371 | _T_108; // @[Decode.scala 15:30]
  assign _T_373 = _T_372 | _T_110; // @[Decode.scala 15:30]
  assign _T_374 = _T_373 | _T_112; // @[Decode.scala 15:30]
  assign _T_375 = _T_374 | _T_114; // @[Decode.scala 15:30]
  assign _T_376 = _T_375 | _T_116; // @[Decode.scala 15:30]
  assign _T_377 = _T_376 | _T_118; // @[Decode.scala 15:30]
  assign _T_378 = _T_377 | _T_120; // @[Decode.scala 15:30]
  assign _T_379 = _T_378 | _T_122; // @[Decode.scala 15:30]
  assign _T_380 = _T_379 | _T_124; // @[Decode.scala 15:30]
  assign _T_381 = _T_380 | _T_126; // @[Decode.scala 15:30]
  assign _T_382 = _T_381 | _T_128; // @[Decode.scala 15:30]
  assign _T_383 = _T_382 | _T_130; // @[Decode.scala 15:30]
  assign _T_384 = _T_383 | _T_132; // @[Decode.scala 15:30]
  assign _T_385 = _T_384 | _T_134; // @[Decode.scala 15:30]
  assign _T_386 = _T_385 | _T_136; // @[Decode.scala 15:30]
  assign _T_387 = _T_386 | _T_138; // @[Decode.scala 15:30]
  assign _T_388 = _T_387 | _T_140; // @[Decode.scala 15:30]
  assign _T_389 = _T_388 | _T_142; // @[Decode.scala 15:30]
  assign _T_390 = _T_389 | _T_144; // @[Decode.scala 15:30]
  assign _T_391 = _T_390 | _T_146; // @[Decode.scala 15:30]
  assign _T_392 = _T_391 | _T_148; // @[Decode.scala 15:30]
  assign _T_393 = _T_392 | _T_150; // @[Decode.scala 15:30]
  assign _T_394 = _T_393 | _T_152; // @[Decode.scala 15:30]
  assign _T_395 = _T_394 | _T_154; // @[Decode.scala 15:30]
  assign _T_396 = _T_395 | _T_156; // @[Decode.scala 15:30]
  assign _T_397 = _T_396 | _T_158; // @[Decode.scala 15:30]
  assign _T_398 = _T_397 | _T_160; // @[Decode.scala 15:30]
  assign _T_399 = _T_398 | _T_162; // @[Decode.scala 15:30]
  assign _T_400 = _T_399 | _T_164; // @[Decode.scala 15:30]
  assign _T_401 = _T_400 | _T_166; // @[Decode.scala 15:30]
  assign _T_402 = _T_401 | _T_168; // @[Decode.scala 15:30]
  assign _T_403 = _T_402 | _T_170; // @[Decode.scala 15:30]
  assign _T_404 = _T_403 | _T_172; // @[Decode.scala 15:30]
  assign _T_405 = _T_404 | _T_174; // @[Decode.scala 15:30]
  assign _T_406 = _T_405 | _T_176; // @[Decode.scala 15:30]
  assign _T_407 = _T_406 | _T_178; // @[Decode.scala 15:30]
  assign _T_408 = _T_407 | _T_180; // @[Decode.scala 15:30]
  assign _T_409 = _T_408 | _T_182; // @[Decode.scala 15:30]
  assign _T_410 = _T_409 | _T_184; // @[Decode.scala 15:30]
  assign _T_411 = _T_410 | _T_186; // @[Decode.scala 15:30]
  assign _T_412 = _T_411 | _T_188; // @[Decode.scala 15:30]
  assign _T_413 = _T_412 | _T_190; // @[Decode.scala 15:30]
  assign _T_414 = _T_413 | _T_192; // @[Decode.scala 15:30]
  assign _T_415 = _T_414 | _T_194; // @[Decode.scala 15:30]
  assign _T_416 = _T_415 | _T_196; // @[Decode.scala 15:30]
  assign _T_417 = _T_416 | _T_198; // @[Decode.scala 15:30]
  assign _T_418 = _T_417 | _T_200; // @[Decode.scala 15:30]
  assign _T_419 = _T_418 | _T_202; // @[Decode.scala 15:30]
  assign _T_420 = _T_419 | _T_204; // @[Decode.scala 15:30]
  assign _T_421 = _T_420 | _T_206; // @[Decode.scala 15:30]
  assign _T_422 = _T_421 | _T_208; // @[Decode.scala 15:30]
  assign _T_423 = _T_422 | _T_210; // @[Decode.scala 15:30]
  assign _T_424 = _T_423 | _T_212; // @[Decode.scala 15:30]
  assign _T_425 = _T_424 | _T_214; // @[Decode.scala 15:30]
  assign _T_426 = _T_425 | _T_216; // @[Decode.scala 15:30]
  assign _T_427 = _T_426 | _T_218; // @[Decode.scala 15:30]
  assign _T_428 = _T_427 | _T_220; // @[Decode.scala 15:30]
  assign _T_429 = _T_428 | _T_222; // @[Decode.scala 15:30]
  assign _T_430 = _T_429 | _T_224; // @[Decode.scala 15:30]
  assign _T_431 = _T_430 | _T_226; // @[Decode.scala 15:30]
  assign _T_432 = _T_431 | _T_228; // @[Decode.scala 15:30]
  assign _T_433 = _T_432 | _T_229; // @[Decode.scala 15:30]
  assign _T_434 = _T_433 | _T_230; // @[Decode.scala 15:30]
  assign _T_435 = _T_434 | _T_232; // @[Decode.scala 15:30]
  assign _T_436 = _T_435 | _T_234; // @[Decode.scala 15:30]
  assign _T_437 = _T_436 | _T_236; // @[Decode.scala 15:30]
  assign _T_438 = _T_437 | _T_238; // @[Decode.scala 15:30]
  assign _T_439 = _T_438 | _T_240; // @[Decode.scala 15:30]
  assign _T_440 = _T_439 | _T_242; // @[Decode.scala 15:30]
  assign _T_441 = _T_440 | _T_244; // @[Decode.scala 15:30]
  assign _T_442 = _T_441 | _T_246; // @[Decode.scala 15:30]
  assign _T_443 = _T_442 | _T_248; // @[Decode.scala 15:30]
  assign _T_444 = _T_443 | _T_250; // @[Decode.scala 15:30]
  assign _T_445 = _T_444 | _T_252; // @[Decode.scala 15:30]
  assign _T_446 = _T_445 | _T_254; // @[Decode.scala 15:30]
  assign _T_447 = _T_446 | _T_256; // @[Decode.scala 15:30]
  assign _T_448 = _T_447 | _T_258; // @[Decode.scala 15:30]
  assign _T_449 = _T_448 | _T_260; // @[Decode.scala 15:30]
  assign _T_450 = _T_449 | _T_262; // @[Decode.scala 15:30]
  assign _T_451 = _T_450 | _T_264; // @[Decode.scala 15:30]
  assign _T_452 = _T_451 | _T_266; // @[Decode.scala 15:30]
  assign _T_453 = _T_452 | _T_268; // @[Decode.scala 15:30]
  assign _T_454 = _T_453 | _T_270; // @[Decode.scala 15:30]
  assign _T_455 = _T_454 | _T_272; // @[Decode.scala 15:30]
  assign _T_456 = _T_455 | _T_274; // @[Decode.scala 15:30]
  assign _T_457 = _T_456 | _T_276; // @[Decode.scala 15:30]
  assign _T_458 = _T_457 | _T_278; // @[Decode.scala 15:30]
  assign _T_459 = _T_458 | _T_280; // @[Decode.scala 15:30]
  assign _T_460 = _T_459 | _T_282; // @[Decode.scala 15:30]
  assign _T_461 = _T_460 | _T_284; // @[Decode.scala 15:30]
  assign _T_462 = _T_461 | _T_286; // @[Decode.scala 15:30]
  assign _T_463 = _T_462 | _T_288; // @[Decode.scala 15:30]
  assign _T_464 = _T_463 | _T_290; // @[Decode.scala 15:30]
  assign _T_465 = _T_464 | _T_292; // @[Decode.scala 15:30]
  assign _T_466 = _T_465 | _T_294; // @[Decode.scala 15:30]
  assign _T_467 = _T_466 | _T_296; // @[Decode.scala 15:30]
  assign _T_468 = _T_467 | _T_298; // @[Decode.scala 15:30]
  assign _T_469 = _T_468 | _T_300; // @[Decode.scala 15:30]
  assign _T_470 = _T_469 | _T_302; // @[Decode.scala 15:30]
  assign _T_471 = _T_470 | _T_303; // @[Decode.scala 15:30]
  assign _T_472 = _T_471 | _T_304; // @[Decode.scala 15:30]
  assign _T_473 = _T_472 | _T_305; // @[Decode.scala 15:30]
  assign _T_474 = _T_473 | _T_306; // @[Decode.scala 15:30]
  assign _T_475 = _T_474 | _T_307; // @[Decode.scala 15:30]
  assign _T_476 = _T_475 | _T_309; // @[Decode.scala 15:30]
  assign _T_477 = _T_476 | _T_311; // @[Decode.scala 15:30]
  assign _T_478 = _T_477 | _T_313; // @[Decode.scala 15:30]
  assign _T_479 = _T_478 | _T_315; // @[Decode.scala 15:30]
  assign _T_480 = _T_479 | _T_317; // @[Decode.scala 15:30]
  assign id_ctrl_legal = _T_480 | _T_319; // @[Decode.scala 15:30]
  assign _T_482 = ibuf_io_inst_0_bits_inst_bits & 32'h5c; // @[Decode.scala 14:65]
  assign _T_483 = _T_482 == 32'h4; // @[Decode.scala 14:121]
  assign _T_484 = ibuf_io_inst_0_bits_inst_bits & 32'h60; // @[Decode.scala 14:65]
  assign _T_485 = _T_484 == 32'h40; // @[Decode.scala 14:121]
  assign id_ctrl_fp = _T_483 | _T_485; // @[Decode.scala 15:30]
  assign _T_488 = ibuf_io_inst_0_bits_inst_bits & 32'h74; // @[Decode.scala 14:65]
  assign id_ctrl_branch = _T_488 == 32'h60; // @[Decode.scala 14:121]
  assign _T_491 = ibuf_io_inst_0_bits_inst_bits & 32'h68; // @[Decode.scala 14:65]
  assign id_ctrl_jal = _T_491 == 32'h68; // @[Decode.scala 14:121]
  assign _T_494 = ibuf_io_inst_0_bits_inst_bits & 32'h203c; // @[Decode.scala 14:65]
  assign id_ctrl_jalr = _T_494 == 32'h24; // @[Decode.scala 14:121]
  assign _T_497 = ibuf_io_inst_0_bits_inst_bits & 32'h64; // @[Decode.scala 14:65]
  assign _T_498 = _T_497 == 32'h20; // @[Decode.scala 14:121]
  assign _T_499 = ibuf_io_inst_0_bits_inst_bits & 32'h34; // @[Decode.scala 14:65]
  assign _T_500 = _T_499 == 32'h20; // @[Decode.scala 14:121]
  assign _T_501 = ibuf_io_inst_0_bits_inst_bits & 32'h2048; // @[Decode.scala 14:65]
  assign _T_502 = _T_501 == 32'h2008; // @[Decode.scala 14:121]
  assign _T_503 = ibuf_io_inst_0_bits_inst_bits & 32'h42003024; // @[Decode.scala 14:65]
  assign _T_504 = _T_503 == 32'h2000020; // @[Decode.scala 14:121]
  assign _T_506 = _T_498 | _T_500; // @[Decode.scala 15:30]
  assign _T_507 = _T_506 | _T_502; // @[Decode.scala 15:30]
  assign id_ctrl_rxs2 = _T_507 | _T_504; // @[Decode.scala 15:30]
  assign _T_509 = ibuf_io_inst_0_bits_inst_bits & 32'h44; // @[Decode.scala 14:65]
  assign _T_510 = _T_509 == 32'h0; // @[Decode.scala 14:121]
  assign _T_511 = ibuf_io_inst_0_bits_inst_bits & 32'h4024; // @[Decode.scala 14:65]
  assign _T_512 = _T_511 == 32'h20; // @[Decode.scala 14:121]
  assign _T_513 = ibuf_io_inst_0_bits_inst_bits & 32'h38; // @[Decode.scala 14:65]
  assign _T_514 = _T_513 == 32'h20; // @[Decode.scala 14:121]
  assign _T_515 = ibuf_io_inst_0_bits_inst_bits & 32'h2050; // @[Decode.scala 14:65]
  assign _T_516 = _T_515 == 32'h2000; // @[Decode.scala 14:121]
  assign _T_517 = ibuf_io_inst_0_bits_inst_bits & 32'h90000034; // @[Decode.scala 14:65]
  assign _T_518 = _T_517 == 32'h90000010; // @[Decode.scala 14:121]
  assign _T_520 = _T_510 | _T_512; // @[Decode.scala 15:30]
  assign _T_521 = _T_520 | _T_514; // @[Decode.scala 15:30]
  assign _T_522 = _T_521 | _T_516; // @[Decode.scala 15:30]
  assign id_ctrl_rxs1 = _T_522 | _T_518; // @[Decode.scala 15:30]
  assign _T_524 = ibuf_io_inst_0_bits_inst_bits & 32'h58; // @[Decode.scala 14:65]
  assign _T_525 = _T_524 == 32'h0; // @[Decode.scala 14:121]
  assign _T_526 = ibuf_io_inst_0_bits_inst_bits & 32'h20; // @[Decode.scala 14:65]
  assign _T_527 = _T_526 == 32'h0; // @[Decode.scala 14:121]
  assign _T_528 = ibuf_io_inst_0_bits_inst_bits & 32'hc; // @[Decode.scala 14:65]
  assign _T_529 = _T_528 == 32'h4; // @[Decode.scala 14:121]
  assign _T_530 = ibuf_io_inst_0_bits_inst_bits & 32'h48; // @[Decode.scala 14:65]
  assign _T_531 = _T_530 == 32'h48; // @[Decode.scala 14:121]
  assign _T_532 = ibuf_io_inst_0_bits_inst_bits & 32'h4050; // @[Decode.scala 14:65]
  assign _T_533 = _T_532 == 32'h4050; // @[Decode.scala 14:121]
  assign _T_535 = _T_525 | _T_527; // @[Decode.scala 15:30]
  assign _T_536 = _T_535 | _T_529; // @[Decode.scala 15:30]
  assign _T_537 = _T_536 | _T_531; // @[Decode.scala 15:30]
  assign _T_538 = _T_537 | _T_533; // @[Decode.scala 15:30]
  assign _T_540 = _T_530 == 32'h0; // @[Decode.scala 14:121]
  assign _T_541 = ibuf_io_inst_0_bits_inst_bits & 32'h18; // @[Decode.scala 14:65]
  assign _T_542 = _T_541 == 32'h0; // @[Decode.scala 14:121]
  assign _T_543 = ibuf_io_inst_0_bits_inst_bits & 32'h4008; // @[Decode.scala 14:65]
  assign _T_544 = _T_543 == 32'h4000; // @[Decode.scala 14:121]
  assign _T_546 = _T_540 | _T_510; // @[Decode.scala 15:30]
  assign _T_547 = _T_546 | _T_542; // @[Decode.scala 15:30]
  assign _T_548 = _T_547 | _T_544; // @[Decode.scala 15:30]
  assign id_ctrl_sel_alu2 = {_T_548,_T_538}; // @[Cat.scala 29:58]
  assign _T_550 = ibuf_io_inst_0_bits_inst_bits & 32'h4004; // @[Decode.scala 14:65]
  assign _T_551 = _T_550 == 32'h0; // @[Decode.scala 14:121]
  assign _T_552 = ibuf_io_inst_0_bits_inst_bits & 32'h50; // @[Decode.scala 14:65]
  assign _T_553 = _T_552 == 32'h0; // @[Decode.scala 14:121]
  assign _T_554 = ibuf_io_inst_0_bits_inst_bits & 32'h24; // @[Decode.scala 14:65]
  assign _T_555 = _T_554 == 32'h0; // @[Decode.scala 14:121]
  assign _T_557 = _T_551 | _T_553; // @[Decode.scala 15:30]
  assign _T_558 = _T_557 | _T_510; // @[Decode.scala 15:30]
  assign _T_559 = _T_558 | _T_555; // @[Decode.scala 15:30]
  assign _T_560 = _T_559 | _T_542; // @[Decode.scala 15:30]
  assign _T_562 = _T_499 == 32'h14; // @[Decode.scala 14:121]
  assign _T_564 = _T_562 | _T_531; // @[Decode.scala 15:30]
  assign id_ctrl_sel_alu1 = {_T_564,_T_560}; // @[Cat.scala 29:58]
  assign _T_567 = _T_541 == 32'h8; // @[Decode.scala 14:121]
  assign _T_569 = _T_509 == 32'h40; // @[Decode.scala 14:121]
  assign _T_571 = _T_567 | _T_569; // @[Decode.scala 15:30]
  assign _T_572 = ibuf_io_inst_0_bits_inst_bits & 32'h14; // @[Decode.scala 14:65]
  assign _T_573 = _T_572 == 32'h14; // @[Decode.scala 14:121]
  assign _T_575 = _T_567 | _T_573; // @[Decode.scala 15:30]
  assign _T_576 = ibuf_io_inst_0_bits_inst_bits & 32'h30; // @[Decode.scala 14:65]
  assign _T_577 = _T_576 == 32'h0; // @[Decode.scala 14:121]
  assign _T_578 = ibuf_io_inst_0_bits_inst_bits & 32'h201c; // @[Decode.scala 14:65]
  assign _T_579 = _T_578 == 32'h4; // @[Decode.scala 14:121]
  assign _T_581 = _T_572 == 32'h10; // @[Decode.scala 14:121]
  assign _T_583 = _T_577 | _T_579; // @[Decode.scala 15:30]
  assign _T_584 = _T_583 | _T_581; // @[Decode.scala 15:30]
  assign id_ctrl_sel_imm = {_T_584,_T_575,_T_571}; // @[Cat.scala 29:58]
  assign _T_587 = ibuf_io_inst_0_bits_inst_bits & 32'h10; // @[Decode.scala 14:65]
  assign _T_588 = _T_587 == 32'h0; // @[Decode.scala 14:121]
  assign _T_589 = ibuf_io_inst_0_bits_inst_bits & 32'h8; // @[Decode.scala 14:65]
  assign _T_590 = _T_589 == 32'h0; // @[Decode.scala 14:121]
  assign id_ctrl_alu_dw = _T_588 | _T_590; // @[Decode.scala 15:30]
  assign _T_593 = ibuf_io_inst_0_bits_inst_bits & 32'h3054; // @[Decode.scala 14:65]
  assign _T_594 = _T_593 == 32'h1010; // @[Decode.scala 14:121]
  assign _T_595 = ibuf_io_inst_0_bits_inst_bits & 32'h1058; // @[Decode.scala 14:65]
  assign _T_596 = _T_595 == 32'h1040; // @[Decode.scala 14:121]
  assign _T_597 = ibuf_io_inst_0_bits_inst_bits & 32'h7044; // @[Decode.scala 14:65]
  assign _T_598 = _T_597 == 32'h7000; // @[Decode.scala 14:121]
  assign _T_599 = ibuf_io_inst_0_bits_inst_bits & 32'h2001074; // @[Decode.scala 14:65]
  assign _T_600 = _T_599 == 32'h2001030; // @[Decode.scala 14:121]
  assign _T_602 = _T_594 | _T_596; // @[Decode.scala 15:30]
  assign _T_603 = _T_602 | _T_598; // @[Decode.scala 15:30]
  assign _T_604 = _T_603 | _T_600; // @[Decode.scala 15:30]
  assign _T_605 = ibuf_io_inst_0_bits_inst_bits & 32'h4054; // @[Decode.scala 14:65]
  assign _T_606 = _T_605 == 32'h40; // @[Decode.scala 14:121]
  assign _T_607 = ibuf_io_inst_0_bits_inst_bits & 32'h2058; // @[Decode.scala 14:65]
  assign _T_608 = _T_607 == 32'h2040; // @[Decode.scala 14:121]
  assign _T_610 = _T_593 == 32'h3010; // @[Decode.scala 14:121]
  assign _T_611 = ibuf_io_inst_0_bits_inst_bits & 32'h6054; // @[Decode.scala 14:65]
  assign _T_612 = _T_611 == 32'h6010; // @[Decode.scala 14:121]
  assign _T_613 = ibuf_io_inst_0_bits_inst_bits & 32'h2002074; // @[Decode.scala 14:65]
  assign _T_614 = _T_613 == 32'h2002030; // @[Decode.scala 14:121]
  assign _T_615 = ibuf_io_inst_0_bits_inst_bits & 32'h40003034; // @[Decode.scala 14:65]
  assign _T_616 = _T_615 == 32'h40000030; // @[Decode.scala 14:121]
  assign _T_617 = ibuf_io_inst_0_bits_inst_bits & 32'h40001054; // @[Decode.scala 14:65]
  assign _T_618 = _T_617 == 32'h40001010; // @[Decode.scala 14:121]
  assign _T_620 = _T_606 | _T_608; // @[Decode.scala 15:30]
  assign _T_621 = _T_620 | _T_610; // @[Decode.scala 15:30]
  assign _T_622 = _T_621 | _T_612; // @[Decode.scala 15:30]
  assign _T_623 = _T_622 | _T_614; // @[Decode.scala 15:30]
  assign _T_624 = _T_623 | _T_616; // @[Decode.scala 15:30]
  assign _T_625 = _T_624 | _T_618; // @[Decode.scala 15:30]
  assign _T_626 = ibuf_io_inst_0_bits_inst_bits & 32'h2002054; // @[Decode.scala 14:65]
  assign _T_627 = _T_626 == 32'h2010; // @[Decode.scala 14:121]
  assign _T_628 = ibuf_io_inst_0_bits_inst_bits & 32'h2034; // @[Decode.scala 14:65]
  assign _T_629 = _T_628 == 32'h2010; // @[Decode.scala 14:121]
  assign _T_630 = ibuf_io_inst_0_bits_inst_bits & 32'h40004054; // @[Decode.scala 14:65]
  assign _T_631 = _T_630 == 32'h4010; // @[Decode.scala 14:121]
  assign _T_632 = ibuf_io_inst_0_bits_inst_bits & 32'h5054; // @[Decode.scala 14:65]
  assign _T_633 = _T_632 == 32'h4010; // @[Decode.scala 14:121]
  assign _T_634 = ibuf_io_inst_0_bits_inst_bits & 32'h4058; // @[Decode.scala 14:65]
  assign _T_635 = _T_634 == 32'h4040; // @[Decode.scala 14:121]
  assign _T_637 = _T_627 | _T_629; // @[Decode.scala 15:30]
  assign _T_638 = _T_637 | _T_631; // @[Decode.scala 15:30]
  assign _T_639 = _T_638 | _T_633; // @[Decode.scala 15:30]
  assign _T_640 = _T_639 | _T_635; // @[Decode.scala 15:30]
  assign _T_641 = ibuf_io_inst_0_bits_inst_bits & 32'h2006054; // @[Decode.scala 14:65]
  assign _T_642 = _T_641 == 32'h2010; // @[Decode.scala 14:121]
  assign _T_643 = ibuf_io_inst_0_bits_inst_bits & 32'h6034; // @[Decode.scala 14:65]
  assign _T_644 = _T_643 == 32'h2010; // @[Decode.scala 14:121]
  assign _T_645 = ibuf_io_inst_0_bits_inst_bits & 32'h40003054; // @[Decode.scala 14:65]
  assign _T_646 = _T_645 == 32'h40001010; // @[Decode.scala 14:121]
  assign _T_648 = _T_642 | _T_644; // @[Decode.scala 15:30]
  assign _T_649 = _T_648 | _T_635; // @[Decode.scala 15:30]
  assign _T_650 = _T_649 | _T_616; // @[Decode.scala 15:30]
  assign _T_651 = _T_650 | _T_646; // @[Decode.scala 15:30]
  assign id_ctrl_alu_fn = {_T_651,_T_640,_T_625,_T_604}; // @[Cat.scala 29:58]
  assign _T_656 = _T_30 | _T_32; // @[Decode.scala 15:30]
  assign _T_657 = _T_656 | _T_34; // @[Decode.scala 15:30]
  assign _T_658 = _T_657 | _T_36; // @[Decode.scala 15:30]
  assign _T_659 = _T_658 | _T_38; // @[Decode.scala 15:30]
  assign _T_660 = _T_659 | _T_40; // @[Decode.scala 15:30]
  assign _T_661 = _T_660 | _T_42; // @[Decode.scala 15:30]
  assign _T_662 = _T_661 | _T_44; // @[Decode.scala 15:30]
  assign _T_663 = _T_662 | _T_46; // @[Decode.scala 15:30]
  assign _T_664 = _T_663 | _T_48; // @[Decode.scala 15:30]
  assign _T_665 = _T_664 | _T_50; // @[Decode.scala 15:30]
  assign _T_666 = _T_665 | _T_52; // @[Decode.scala 15:30]
  assign _T_667 = _T_666 | _T_54; // @[Decode.scala 15:30]
  assign _T_668 = _T_667 | _T_56; // @[Decode.scala 15:30]
  assign _T_669 = _T_668 | _T_58; // @[Decode.scala 15:30]
  assign _T_670 = _T_669 | _T_60; // @[Decode.scala 15:30]
  assign _T_671 = _T_670 | _T_62; // @[Decode.scala 15:30]
  assign _T_672 = _T_671 | _T_64; // @[Decode.scala 15:30]
  assign _T_673 = _T_672 | _T_66; // @[Decode.scala 15:30]
  assign _T_674 = _T_673 | _T_68; // @[Decode.scala 15:30]
  assign _T_675 = _T_674 | _T_70; // @[Decode.scala 15:30]
  assign _T_676 = _T_675 | _T_72; // @[Decode.scala 15:30]
  assign _T_677 = _T_676 | _T_118; // @[Decode.scala 15:30]
  assign _T_678 = _T_677 | _T_120; // @[Decode.scala 15:30]
  assign _T_679 = _T_678 | _T_178; // @[Decode.scala 15:30]
  assign _T_680 = _T_679 | _T_180; // @[Decode.scala 15:30]
  assign _T_681 = _T_680 | _T_198; // @[Decode.scala 15:30]
  assign _T_682 = _T_681 | _T_200; // @[Decode.scala 15:30]
  assign _T_683 = _T_682 | _T_202; // @[Decode.scala 15:30]
  assign _T_684 = _T_683 | _T_228; // @[Decode.scala 15:30]
  assign _T_685 = _T_684 | _T_252; // @[Decode.scala 15:30]
  assign _T_686 = _T_685 | _T_254; // @[Decode.scala 15:30]
  assign _T_687 = _T_686 | _T_256; // @[Decode.scala 15:30]
  assign _T_688 = _T_687 | _T_258; // @[Decode.scala 15:30]
  assign _T_689 = _T_688 | _T_260; // @[Decode.scala 15:30]
  assign _T_690 = _T_689 | _T_262; // @[Decode.scala 15:30]
  assign _T_691 = _T_690 | _T_264; // @[Decode.scala 15:30]
  assign id_ctrl_mem = _T_691 | _T_266; // @[Decode.scala 15:30]
  assign _T_694 = _T_491 == 32'h20; // @[Decode.scala 14:121]
  assign _T_695 = ibuf_io_inst_0_bits_inst_bits & 32'h18000020; // @[Decode.scala 14:65]
  assign _T_696 = _T_695 == 32'h18000020; // @[Decode.scala 14:121]
  assign _T_697 = ibuf_io_inst_0_bits_inst_bits & 32'h20000020; // @[Decode.scala 14:65]
  assign _T_698 = _T_697 == 32'h20000020; // @[Decode.scala 14:121]
  assign _T_700 = _T_694 | _T_696; // @[Decode.scala 15:30]
  assign _T_701 = _T_700 | _T_698; // @[Decode.scala 15:30]
  assign _T_702 = ibuf_io_inst_0_bits_inst_bits & 32'h10000008; // @[Decode.scala 14:65]
  assign _T_703 = _T_702 == 32'h10000008; // @[Decode.scala 14:121]
  assign _T_704 = ibuf_io_inst_0_bits_inst_bits & 32'h40000008; // @[Decode.scala 14:65]
  assign _T_705 = _T_704 == 32'h40000008; // @[Decode.scala 14:121]
  assign _T_707 = _T_703 | _T_705; // @[Decode.scala 15:30]
  assign _T_708 = ibuf_io_inst_0_bits_inst_bits & 32'h40; // @[Decode.scala 14:65]
  assign _T_709 = _T_708 == 32'h40; // @[Decode.scala 14:121]
  assign _T_710 = ibuf_io_inst_0_bits_inst_bits & 32'h8000008; // @[Decode.scala 14:65]
  assign _T_711 = _T_710 == 32'h8000008; // @[Decode.scala 14:121]
  assign _T_712 = ibuf_io_inst_0_bits_inst_bits & 32'h80000008; // @[Decode.scala 14:65]
  assign _T_713 = _T_712 == 32'h80000008; // @[Decode.scala 14:121]
  assign _T_715 = _T_709 | _T_711; // @[Decode.scala 15:30]
  assign _T_716 = _T_715 | _T_703; // @[Decode.scala 15:30]
  assign _T_717 = _T_716 | _T_713; // @[Decode.scala 15:30]
  assign _T_718 = ibuf_io_inst_0_bits_inst_bits & 32'h18000008; // @[Decode.scala 14:65]
  assign _T_719 = _T_718 == 32'h8; // @[Decode.scala 14:121]
  assign id_ctrl_mem_cmd = {_T_709,_T_719,_T_717,_T_707,_T_701}; // @[Cat.scala 29:58]
  assign _T_726 = ibuf_io_inst_0_bits_inst_bits & 32'h80000060; // @[Decode.scala 14:65]
  assign _T_727 = _T_726 == 32'h40; // @[Decode.scala 14:121]
  assign _T_728 = ibuf_io_inst_0_bits_inst_bits & 32'h10000060; // @[Decode.scala 14:65]
  assign _T_729 = _T_728 == 32'h40; // @[Decode.scala 14:121]
  assign _T_730 = ibuf_io_inst_0_bits_inst_bits & 32'h70; // @[Decode.scala 14:65]
  assign id_ctrl_rfs3 = _T_730 == 32'h40; // @[Decode.scala 14:121]
  assign _T_733 = _T_727 | _T_729; // @[Decode.scala 15:30]
  assign id_ctrl_rfs1 = _T_733 | id_ctrl_rfs3; // @[Decode.scala 15:30]
  assign _T_735 = ibuf_io_inst_0_bits_inst_bits & 32'h7c; // @[Decode.scala 14:65]
  assign _T_736 = _T_735 == 32'h24; // @[Decode.scala 14:121]
  assign _T_737 = ibuf_io_inst_0_bits_inst_bits & 32'h40000060; // @[Decode.scala 14:65]
  assign _T_738 = _T_737 == 32'h40; // @[Decode.scala 14:121]
  assign _T_739 = ibuf_io_inst_0_bits_inst_bits & 32'h90000060; // @[Decode.scala 14:65]
  assign _T_740 = _T_739 == 32'h10000040; // @[Decode.scala 14:121]
  assign _T_742 = _T_736 | _T_738; // @[Decode.scala 15:30]
  assign _T_743 = _T_742 | id_ctrl_rfs3; // @[Decode.scala 15:30]
  assign id_ctrl_rfs2 = _T_743 | _T_740; // @[Decode.scala 15:30]
  assign _T_746 = ibuf_io_inst_0_bits_inst_bits & 32'h3c; // @[Decode.scala 14:65]
  assign _T_747 = _T_746 == 32'h4; // @[Decode.scala 14:121]
  assign _T_749 = _T_728 == 32'h10000040; // @[Decode.scala 14:121]
  assign _T_751 = _T_747 | _T_727; // @[Decode.scala 15:30]
  assign _T_752 = _T_751 | id_ctrl_rfs3; // @[Decode.scala 15:30]
  assign id_ctrl_wfd = _T_752 | _T_749; // @[Decode.scala 15:30]
  assign _T_754 = ibuf_io_inst_0_bits_inst_bits & 32'h2000074; // @[Decode.scala 14:65]
  assign id_ctrl_div = _T_754 == 32'h2000030; // @[Decode.scala 14:121]
  assign _T_758 = _T_497 == 32'h0; // @[Decode.scala 14:121]
  assign _T_760 = _T_552 == 32'h10; // @[Decode.scala 14:121]
  assign _T_761 = ibuf_io_inst_0_bits_inst_bits & 32'h2024; // @[Decode.scala 14:65]
  assign _T_762 = _T_761 == 32'h24; // @[Decode.scala 14:121]
  assign _T_763 = ibuf_io_inst_0_bits_inst_bits & 32'h28; // @[Decode.scala 14:65]
  assign _T_764 = _T_763 == 32'h28; // @[Decode.scala 14:121]
  assign _T_765 = ibuf_io_inst_0_bits_inst_bits & 32'h1030; // @[Decode.scala 14:65]
  assign _T_766 = _T_765 == 32'h1030; // @[Decode.scala 14:121]
  assign _T_767 = ibuf_io_inst_0_bits_inst_bits & 32'h2030; // @[Decode.scala 14:65]
  assign _T_768 = _T_767 == 32'h2030; // @[Decode.scala 14:121]
  assign _T_769 = ibuf_io_inst_0_bits_inst_bits & 32'h90000010; // @[Decode.scala 14:65]
  assign _T_770 = _T_769 == 32'h80000010; // @[Decode.scala 14:121]
  assign _T_772 = _T_758 | _T_760; // @[Decode.scala 15:30]
  assign _T_773 = _T_772 | _T_762; // @[Decode.scala 15:30]
  assign _T_774 = _T_773 | _T_764; // @[Decode.scala 15:30]
  assign _T_775 = _T_774 | _T_766; // @[Decode.scala 15:30]
  assign _T_776 = _T_775 | _T_768; // @[Decode.scala 15:30]
  assign id_ctrl_wxd = _T_776 | _T_770; // @[Decode.scala 15:30]
  assign _T_778 = ibuf_io_inst_0_bits_inst_bits & 32'h1070; // @[Decode.scala 14:65]
  assign _T_779 = _T_778 == 32'h1070; // @[Decode.scala 14:121]
  assign _T_781 = ibuf_io_inst_0_bits_inst_bits & 32'h2070; // @[Decode.scala 14:65]
  assign _T_782 = _T_781 == 32'h2070; // @[Decode.scala 14:121]
  assign _T_784 = ibuf_io_inst_0_bits_inst_bits & 32'h10000070; // @[Decode.scala 14:65]
  assign _T_785 = _T_784 == 32'h70; // @[Decode.scala 14:121]
  assign _T_786 = ibuf_io_inst_0_bits_inst_bits & 32'h12000034; // @[Decode.scala 14:65]
  assign _T_787 = _T_786 == 32'h10000030; // @[Decode.scala 14:121]
  assign _T_788 = ibuf_io_inst_0_bits_inst_bits & 32'he0000050; // @[Decode.scala 14:65]
  assign _T_789 = _T_788 == 32'h60000050; // @[Decode.scala 14:121]
  assign _T_791 = _T_785 | _T_779; // @[Decode.scala 15:30]
  assign _T_792 = _T_791 | _T_782; // @[Decode.scala 15:30]
  assign _T_793 = _T_792 | _T_787; // @[Decode.scala 15:30]
  assign _T_794 = _T_793 | _T_789; // @[Decode.scala 15:30]
  assign id_ctrl_csr = {_T_794,_T_782,_T_779}; // @[Cat.scala 29:58]
  assign _T_797 = ibuf_io_inst_0_bits_inst_bits & 32'h3058; // @[Decode.scala 14:65]
  assign id_ctrl_fence_i = _T_797 == 32'h1008; // @[Decode.scala 14:121]
  assign id_ctrl_fence = _T_607 == 32'h8; // @[Decode.scala 14:121]
  assign _T_803 = ibuf_io_inst_0_bits_inst_bits & 32'h6048; // @[Decode.scala 14:65]
  assign id_ctrl_amo = _T_803 == 32'h2008; // @[Decode.scala 14:121]
  assign _T_806 = ibuf_io_inst_0_bits_inst_bits & 32'h105c; // @[Decode.scala 14:65]
  assign _T_807 = _T_806 == 32'h1004; // @[Decode.scala 14:121]
  assign _T_808 = ibuf_io_inst_0_bits_inst_bits & 32'h2000060; // @[Decode.scala 14:65]
  assign _T_809 = _T_808 == 32'h2000040; // @[Decode.scala 14:121]
  assign _T_810 = ibuf_io_inst_0_bits_inst_bits & 32'hd0000070; // @[Decode.scala 14:65]
  assign _T_811 = _T_810 == 32'h40000050; // @[Decode.scala 14:121]
  assign _T_813 = _T_807 | _T_809; // @[Decode.scala 15:30]
  assign id_ctrl_dp = _T_813 | _T_811; // @[Decode.scala 15:30]
  assign id_raddr3 = ibuf_io_inst_0_bits_inst_rs3; // @[RocketCore.scala 261:72]
  assign id_raddr2 = ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 261:72]
  assign id_raddr1 = ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 261:72]
  assign id_waddr = ibuf_io_inst_0_bits_inst_rd; // @[RocketCore.scala 261:72]
  assign _T_816 = id_raddr1 == 5'h0; // @[RocketCore.scala 1021:45]
  assign _T_821 = _T_815__T_820_data; // @[RocketCore.scala 1021:25]
  assign _T_827 = _T_815__T_826_data; // @[RocketCore.scala 1021:25]
  assign _T_894 = id_ctrl_csr == 3'h6; // @[package.scala 15:47]
  assign _T_895 = id_ctrl_csr == 3'h7; // @[package.scala 15:47]
  assign _T_896 = id_ctrl_csr == 3'h5; // @[package.scala 15:47]
  assign _T_897 = _T_894 | _T_895; // @[package.scala 64:59]
  assign id_csr_en = _T_897 | _T_896; // @[package.scala 64:59]
  assign id_system_insn = id_ctrl_csr == 3'h4; // @[RocketCore.scala 278:36]
  assign id_csr_ren = _T_897 & _T_816; // @[RocketCore.scala 279:54]
  assign _T_902 = id_ctrl_mem_cmd == 5'h14; // @[RocketCore.scala 281:50]
  assign id_sfence = id_ctrl_mem & _T_902; // @[RocketCore.scala 281:31]
  assign _T_903 = id_sfence | id_system_insn; // @[RocketCore.scala 282:32]
  assign _T_905 = id_csr_en & ~id_csr_ren; // @[RocketCore.scala 282:64]
  assign _T_906 = _T_905 & csr_io_decode_0_write_flush; // @[RocketCore.scala 282:79]
  assign id_csr_flush = _T_903 | _T_906; // @[RocketCore.scala 282:50]
  assign _T_911 = id_ctrl_div & ~csr_io_status_isa[12]; // @[RocketCore.scala 291:34]
  assign _T_912 = ~id_ctrl_legal | _T_911; // @[RocketCore.scala 290:40]
  assign _T_915 = id_ctrl_amo & ~csr_io_status_isa[0]; // @[RocketCore.scala 292:17]
  assign _T_916 = _T_912 | _T_915; // @[RocketCore.scala 291:65]
  assign _T_917 = csr_io_decode_0_fp_illegal | io_fpu_illegal_rm; // @[RocketCore.scala 293:48]
  assign _T_918 = id_ctrl_fp & _T_917; // @[RocketCore.scala 293:16]
  assign _T_919 = _T_916 | _T_918; // @[RocketCore.scala 292:48]
  assign _T_922 = id_ctrl_dp & ~csr_io_status_isa[3]; // @[RocketCore.scala 294:16]
  assign _T_923 = _T_919 | _T_922; // @[RocketCore.scala 293:70]
  assign _T_926 = ibuf_io_inst_0_bits_rvc & ~csr_io_status_isa[2]; // @[RocketCore.scala 295:30]
  assign _T_927 = _T_923 | _T_926; // @[RocketCore.scala 294:47]
  assign _T_947 = ~id_csr_ren & csr_io_decode_0_write_illegal; // @[RocketCore.scala 301:64]
  assign _T_948 = csr_io_decode_0_read_illegal | _T_947; // @[RocketCore.scala 301:49]
  assign _T_949 = id_csr_en & _T_948; // @[RocketCore.scala 301:15]
  assign _T_950 = _T_927 | _T_949; // @[RocketCore.scala 300:81]
  assign _T_953 = _T_903 & csr_io_decode_0_system_illegal; // @[RocketCore.scala 302:65]
  assign _T_954 = ~ibuf_io_inst_0_bits_rvc & _T_953; // @[RocketCore.scala 302:31]
  assign id_illegal_insn = _T_950 | _T_954; // @[RocketCore.scala 301:99]
  assign id_amo_aq = ibuf_io_inst_0_bits_inst_bits[26]; // @[RocketCore.scala 304:29]
  assign id_amo_rl = ibuf_io_inst_0_bits_inst_bits[25]; // @[RocketCore.scala 305:29]
  assign id_fence_succ = ibuf_io_inst_0_bits_inst_bits[23:20]; // @[RocketCore.scala 307:33]
  assign _T_955 = id_ctrl_amo & id_amo_aq; // @[RocketCore.scala 308:52]
  assign id_fence_next = id_ctrl_fence | _T_955; // @[RocketCore.scala 308:37]
  assign id_mem_busy = ~io_dmem_ordered | io_dmem_req_valid; // @[RocketCore.scala 309:38]
  assign _GEN_0 = id_mem_busy ? id_reg_fence : 1'h0; // @[RocketCore.scala 310:23]
  assign _T_965 = id_ctrl_amo & id_amo_rl; // @[RocketCore.scala 315:33]
  assign _T_966 = _T_965 | id_ctrl_fence_i; // @[RocketCore.scala 315:46]
  assign _T_968 = id_reg_fence & id_ctrl_mem; // @[RocketCore.scala 315:81]
  assign _T_969 = _T_966 | _T_968; // @[RocketCore.scala 315:65]
  assign id_do_fence = id_mem_busy & _T_969; // @[RocketCore.scala 315:17]
  assign _T_972 = csr_io_interrupt | bpu_io_debug_if; // @[RocketCore.scala 974:26]
  assign _T_973 = _T_972 | bpu_io_xcpt_if; // @[RocketCore.scala 974:26]
  assign _T_974 = _T_973 | ibuf_io_inst_0_bits_xcpt0_pf_inst; // @[RocketCore.scala 974:26]
  assign _T_975 = _T_974 | ibuf_io_inst_0_bits_xcpt0_ae_inst; // @[RocketCore.scala 974:26]
  assign _T_976 = _T_975 | ibuf_io_inst_0_bits_xcpt1_pf_inst; // @[RocketCore.scala 974:26]
  assign _T_977 = _T_976 | ibuf_io_inst_0_bits_xcpt1_ae_inst; // @[RocketCore.scala 974:26]
  assign id_xcpt = _T_977 | id_illegal_insn; // @[RocketCore.scala 974:26]
  assign _T_978 = ibuf_io_inst_0_bits_xcpt1_ae_inst ? 2'h1 : 2'h2; // @[Mux.scala 47:69]
  assign _T_979 = ibuf_io_inst_0_bits_xcpt1_pf_inst ? 4'hc : {{2'd0}, _T_978}; // @[Mux.scala 47:69]
  assign _T_980 = ibuf_io_inst_0_bits_xcpt0_ae_inst ? 4'h1 : _T_979; // @[Mux.scala 47:69]
  assign _T_981 = ibuf_io_inst_0_bits_xcpt0_pf_inst ? 4'hc : _T_980; // @[Mux.scala 47:69]
  assign _T_982 = bpu_io_xcpt_if ? 4'h3 : _T_981; // @[Mux.scala 47:69]
  assign _T_983 = bpu_io_debug_if ? 4'he : _T_982; // @[Mux.scala 47:69]
  assign ex_waddr = ex_reg_inst[11:7]; // @[RocketCore.scala 351:29]
  assign mem_waddr = mem_reg_inst[11:7]; // @[RocketCore.scala 352:31]
  assign wb_waddr = wb_reg_inst[11:7]; // @[RocketCore.scala 353:29]
  assign _T_997 = ex_reg_valid & ex_ctrl_wxd; // @[RocketCore.scala 356:19]
  assign _T_998 = mem_reg_valid & mem_ctrl_wxd; // @[RocketCore.scala 357:20]
  assign _T_1000 = _T_998 & ~mem_ctrl_mem; // @[RocketCore.scala 357:36]
  assign id_bypass_src_0_0 = 5'h0 == id_raddr1; // @[RocketCore.scala 359:82]
  assign _T_1003 = ex_waddr == id_raddr1; // @[RocketCore.scala 359:82]
  assign id_bypass_src_0_1 = _T_997 & _T_1003; // @[RocketCore.scala 359:74]
  assign _T_1004 = mem_waddr == id_raddr1; // @[RocketCore.scala 359:82]
  assign id_bypass_src_0_2 = _T_1000 & _T_1004; // @[RocketCore.scala 359:74]
  assign id_bypass_src_0_3 = _T_998 & _T_1004; // @[RocketCore.scala 359:74]
  assign id_bypass_src_1_0 = 5'h0 == id_raddr2; // @[RocketCore.scala 359:82]
  assign _T_1007 = ex_waddr == id_raddr2; // @[RocketCore.scala 359:82]
  assign id_bypass_src_1_1 = _T_997 & _T_1007; // @[RocketCore.scala 359:74]
  assign _T_1008 = mem_waddr == id_raddr2; // @[RocketCore.scala 359:82]
  assign id_bypass_src_1_2 = _T_1000 & _T_1008; // @[RocketCore.scala 359:74]
  assign id_bypass_src_1_3 = _T_998 & _T_1008; // @[RocketCore.scala 359:74]
  assign _T_1010 = ex_reg_rs_lsb_0 == 2'h1; // @[package.scala 32:86]
  assign _T_1011 = _T_1010 ? mem_reg_wdata : 64'h0; // @[package.scala 32:76]
  assign _T_1012 = ex_reg_rs_lsb_0 == 2'h2; // @[package.scala 32:86]
  assign _T_1013 = _T_1012 ? wb_reg_wdata : _T_1011; // @[package.scala 32:76]
  assign _T_1014 = ex_reg_rs_lsb_0 == 2'h3; // @[package.scala 32:86]
  assign _T_1015 = _T_1014 ? io_dmem_resp_bits_data_word_bypass : _T_1013; // @[package.scala 32:76]
  assign _T_1016 = {ex_reg_rs_msb_0,ex_reg_rs_lsb_0}; // @[Cat.scala 29:58]
  assign _T_1017 = ex_reg_rs_lsb_1 == 2'h1; // @[package.scala 32:86]
  assign _T_1018 = _T_1017 ? mem_reg_wdata : 64'h0; // @[package.scala 32:76]
  assign _T_1019 = ex_reg_rs_lsb_1 == 2'h2; // @[package.scala 32:86]
  assign _T_1020 = _T_1019 ? wb_reg_wdata : _T_1018; // @[package.scala 32:76]
  assign _T_1021 = ex_reg_rs_lsb_1 == 2'h3; // @[package.scala 32:86]
  assign _T_1022 = _T_1021 ? io_dmem_resp_bits_data_word_bypass : _T_1020; // @[package.scala 32:76]
  assign _T_1023 = {ex_reg_rs_msb_1,ex_reg_rs_lsb_1}; // @[Cat.scala 29:58]
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? _T_1022 : _T_1023; // @[RocketCore.scala 367:14]
  assign _T_1024 = ex_ctrl_sel_imm == 3'h5; // @[RocketCore.scala 1036:24]
  assign _T_1026 = ex_reg_inst[31]; // @[RocketCore.scala 1036:53]
  assign _T_1027 = _T_1024 ? $signed(1'sh0) : $signed(_T_1026); // @[RocketCore.scala 1036:19]
  assign _T_1028 = ex_ctrl_sel_imm == 3'h2; // @[RocketCore.scala 1037:26]
  assign _T_1030 = ex_reg_inst[30:20]; // @[RocketCore.scala 1037:49]
  assign _T_1032 = ex_ctrl_sel_imm != 3'h2; // @[RocketCore.scala 1038:26]
  assign _T_1033 = ex_ctrl_sel_imm != 3'h3; // @[RocketCore.scala 1038:43]
  assign _T_1034 = _T_1032 & _T_1033; // @[RocketCore.scala 1038:36]
  assign _T_1036 = ex_reg_inst[19:12]; // @[RocketCore.scala 1038:73]
  assign _T_1040 = _T_1028 | _T_1024; // @[RocketCore.scala 1039:33]
  assign _T_1041 = ex_ctrl_sel_imm == 3'h3; // @[RocketCore.scala 1040:23]
  assign _T_1043 = ex_reg_inst[20]; // @[RocketCore.scala 1040:44]
  assign _T_1044 = ex_ctrl_sel_imm == 3'h1; // @[RocketCore.scala 1041:23]
  assign _T_1046 = ex_reg_inst[7]; // @[RocketCore.scala 1041:43]
  assign _T_1047 = _T_1044 ? $signed(_T_1046) : $signed(_T_1027); // @[RocketCore.scala 1041:18]
  assign _T_1048 = _T_1041 ? $signed(_T_1043) : $signed(_T_1047); // @[RocketCore.scala 1040:18]
  assign _T_1054 = _T_1040 ? 6'h0 : ex_reg_inst[30:25]; // @[RocketCore.scala 1042:20]
  assign _T_1056 = ex_ctrl_sel_imm == 3'h0; // @[RocketCore.scala 1044:24]
  assign _T_1058 = _T_1056 | _T_1044; // @[RocketCore.scala 1044:34]
  assign _T_1063 = _T_1024 ? ex_reg_inst[19:16] : ex_reg_inst[24:21]; // @[RocketCore.scala 1045:19]
  assign _T_1064 = _T_1058 ? ex_reg_inst[11:8] : _T_1063; // @[RocketCore.scala 1044:19]
  assign _T_1065 = _T_1028 ? 4'h0 : _T_1064; // @[RocketCore.scala 1043:19]
  assign _T_1068 = ex_ctrl_sel_imm == 3'h4; // @[RocketCore.scala 1047:22]
  assign _T_1072 = _T_1024 & ex_reg_inst[15]; // @[RocketCore.scala 1048:17]
  assign _T_1073 = _T_1068 ? ex_reg_inst[20] : _T_1072; // @[RocketCore.scala 1047:17]
  assign _T_1074 = _T_1056 ? ex_reg_inst[7] : _T_1073; // @[RocketCore.scala 1046:17]
  assign _T_1077 = _T_1040 ? $signed(1'sh0) : $signed(_T_1048); // @[Cat.scala 29:58]
  assign _T_1078 = _T_1034 ? $signed({8{_T_1027}}) : $signed(_T_1036); // @[Cat.scala 29:58]
  assign _T_1080 = _T_1028 ? $signed(_T_1030) : $signed({11{_T_1027}}); // @[Cat.scala 29:58]
  assign _T_1081 = _T_1024 ? $signed(1'sh0) : $signed(_T_1026); // @[Cat.scala 29:58]
  assign ex_imm = {_T_1081,_T_1080,_T_1078,_T_1077,_T_1054,_T_1065,_T_1074}; // @[RocketCore.scala 1050:53]
  assign _T_1085 = ex_reg_rs_bypass_0 ? _T_1015 : _T_1016; // @[RocketCore.scala 370:24]
  assign _T_1087 = 2'h1 == ex_ctrl_sel_alu1; // @[Mux.scala 80:60]
  assign _T_1088 = _T_1087 ? $signed(_T_1085) : $signed(64'sh0); // @[Mux.scala 80:57]
  assign _T_1089 = 2'h2 == ex_ctrl_sel_alu1; // @[Mux.scala 80:60]
  assign _T_1090 = ex_reg_rs_bypass_1 ? _T_1022 : _T_1023; // @[RocketCore.scala 373:24]
  assign _T_1091 = ex_reg_rvc ? $signed(4'sh2) : $signed(4'sh4); // @[RocketCore.scala 375:19]
  assign _T_1092 = 2'h2 == ex_ctrl_sel_alu2; // @[Mux.scala 80:60]
  assign _T_1093 = _T_1092 ? $signed(_T_1090) : $signed(64'sh0); // @[Mux.scala 80:57]
  assign _T_1094 = 2'h3 == ex_ctrl_sel_alu2; // @[Mux.scala 80:60]
  assign _T_1095 = _T_1094 ? $signed({{32{ex_imm[31]}},ex_imm}) : $signed(_T_1093); // @[Mux.scala 80:57]
  assign _T_1096 = 2'h1 == ex_ctrl_sel_alu2; // @[Mux.scala 80:60]
  assign _T_1763 = ~ibuf_io_inst_0_valid | ibuf_io_inst_0_bits_replay; // @[RocketCore.scala 776:40]
  assign _T_1764 = _T_1763 | take_pc_mem_wb; // @[RocketCore.scala 776:71]
  assign _T_1568 = id_raddr1 != 5'h0; // @[RocketCore.scala 706:55]
  assign _T_1569 = id_ctrl_rxs1 & _T_1568; // @[RocketCore.scala 706:42]
  assign _T_1616 = id_raddr1 == ex_waddr; // @[RocketCore.scala 726:70]
  assign _T_1617 = _T_1569 & _T_1616; // @[RocketCore.scala 983:27]
  assign _T_1570 = id_raddr2 != 5'h0; // @[RocketCore.scala 707:55]
  assign _T_1571 = id_ctrl_rxs2 & _T_1570; // @[RocketCore.scala 707:42]
  assign _T_1618 = id_raddr2 == ex_waddr; // @[RocketCore.scala 726:70]
  assign _T_1619 = _T_1571 & _T_1618; // @[RocketCore.scala 983:27]
  assign _T_1622 = _T_1617 | _T_1619; // @[RocketCore.scala 983:50]
  assign _T_1572 = id_waddr != 5'h0; // @[RocketCore.scala 708:55]
  assign _T_1573 = id_ctrl_wxd & _T_1572; // @[RocketCore.scala 708:42]
  assign _T_1620 = id_waddr == ex_waddr; // @[RocketCore.scala 726:70]
  assign _T_1621 = _T_1573 & _T_1620; // @[RocketCore.scala 983:27]
  assign _T_1623 = _T_1622 | _T_1621; // @[RocketCore.scala 983:50]
  assign data_hazard_ex = ex_ctrl_wxd & _T_1623; // @[RocketCore.scala 726:36]
  assign _T_1609 = ex_ctrl_csr != 3'h0; // @[RocketCore.scala 725:38]
  assign _T_1610 = _T_1609 | ex_ctrl_jalr; // @[RocketCore.scala 725:48]
  assign _T_1611 = _T_1610 | ex_ctrl_mem; // @[RocketCore.scala 725:64]
  assign _T_1613 = _T_1611 | ex_ctrl_div; // @[RocketCore.scala 725:94]
  assign ex_cannot_bypass = _T_1613 | ex_ctrl_fp; // @[RocketCore.scala 725:109]
  assign _T_1635 = data_hazard_ex & ex_cannot_bypass; // @[RocketCore.scala 728:54]
  assign _T_1625 = io_fpu_dec_ren1 & _T_1616; // @[RocketCore.scala 983:27]
  assign _T_1627 = io_fpu_dec_ren2 & _T_1618; // @[RocketCore.scala 983:27]
  assign _T_1632 = _T_1625 | _T_1627; // @[RocketCore.scala 983:50]
  assign _T_1628 = id_raddr3 == ex_waddr; // @[RocketCore.scala 727:76]
  assign _T_1629 = io_fpu_dec_ren3 & _T_1628; // @[RocketCore.scala 983:27]
  assign _T_1633 = _T_1632 | _T_1629; // @[RocketCore.scala 983:50]
  assign _T_1631 = io_fpu_dec_wen & _T_1620; // @[RocketCore.scala 983:27]
  assign _T_1634 = _T_1633 | _T_1631; // @[RocketCore.scala 983:50]
  assign fp_data_hazard_ex = ex_ctrl_wfd & _T_1634; // @[RocketCore.scala 727:39]
  assign _T_1636 = _T_1635 | fp_data_hazard_ex; // @[RocketCore.scala 728:74]
  assign id_ex_hazard = ex_reg_valid & _T_1636; // @[RocketCore.scala 728:35]
  assign _T_1643 = id_raddr1 == mem_waddr; // @[RocketCore.scala 735:72]
  assign _T_1644 = _T_1569 & _T_1643; // @[RocketCore.scala 983:27]
  assign _T_1645 = id_raddr2 == mem_waddr; // @[RocketCore.scala 735:72]
  assign _T_1646 = _T_1571 & _T_1645; // @[RocketCore.scala 983:27]
  assign _T_1649 = _T_1644 | _T_1646; // @[RocketCore.scala 983:50]
  assign _T_1647 = id_waddr == mem_waddr; // @[RocketCore.scala 735:72]
  assign _T_1648 = _T_1573 & _T_1647; // @[RocketCore.scala 983:27]
  assign _T_1650 = _T_1649 | _T_1648; // @[RocketCore.scala 983:50]
  assign data_hazard_mem = mem_ctrl_wxd & _T_1650; // @[RocketCore.scala 735:38]
  assign _T_1637 = mem_ctrl_csr != 3'h0; // @[RocketCore.scala 734:40]
  assign _T_1638 = mem_ctrl_mem & mem_reg_slow_bypass; // @[RocketCore.scala 734:66]
  assign _T_1639 = _T_1637 | _T_1638; // @[RocketCore.scala 734:50]
  assign _T_1641 = _T_1639 | mem_ctrl_div; // @[RocketCore.scala 734:100]
  assign mem_cannot_bypass = _T_1641 | mem_ctrl_fp; // @[RocketCore.scala 734:116]
  assign _T_1662 = data_hazard_mem & mem_cannot_bypass; // @[RocketCore.scala 737:57]
  assign _T_1652 = io_fpu_dec_ren1 & _T_1643; // @[RocketCore.scala 983:27]
  assign _T_1654 = io_fpu_dec_ren2 & _T_1645; // @[RocketCore.scala 983:27]
  assign _T_1659 = _T_1652 | _T_1654; // @[RocketCore.scala 983:50]
  assign _T_1655 = id_raddr3 == mem_waddr; // @[RocketCore.scala 736:78]
  assign _T_1656 = io_fpu_dec_ren3 & _T_1655; // @[RocketCore.scala 983:27]
  assign _T_1660 = _T_1659 | _T_1656; // @[RocketCore.scala 983:50]
  assign _T_1658 = io_fpu_dec_wen & _T_1647; // @[RocketCore.scala 983:27]
  assign _T_1661 = _T_1660 | _T_1658; // @[RocketCore.scala 983:50]
  assign fp_data_hazard_mem = mem_ctrl_wfd & _T_1661; // @[RocketCore.scala 736:41]
  assign _T_1663 = _T_1662 | fp_data_hazard_mem; // @[RocketCore.scala 737:78]
  assign id_mem_hazard = mem_reg_valid & _T_1663; // @[RocketCore.scala 737:37]
  assign _T_1733 = id_ex_hazard | id_mem_hazard; // @[RocketCore.scala 764:18]
  assign _T_1666 = id_raddr1 == wb_waddr; // @[RocketCore.scala 741:70]
  assign _T_1667 = _T_1569 & _T_1666; // @[RocketCore.scala 983:27]
  assign _T_1668 = id_raddr2 == wb_waddr; // @[RocketCore.scala 741:70]
  assign _T_1669 = _T_1571 & _T_1668; // @[RocketCore.scala 983:27]
  assign _T_1672 = _T_1667 | _T_1669; // @[RocketCore.scala 983:50]
  assign _T_1670 = id_waddr == wb_waddr; // @[RocketCore.scala 741:70]
  assign _T_1671 = _T_1573 & _T_1670; // @[RocketCore.scala 983:27]
  assign _T_1673 = _T_1672 | _T_1671; // @[RocketCore.scala 983:50]
  assign data_hazard_wb = wb_ctrl_wxd & _T_1673; // @[RocketCore.scala 741:36]
  assign wb_dcache_miss = wb_ctrl_mem & ~io_dmem_resp_valid; // @[RocketCore.scala 483:36]
  assign wb_set_sboard = wb_ctrl_div | wb_dcache_miss; // @[RocketCore.scala 628:35]
  assign _T_1685 = data_hazard_wb & wb_set_sboard; // @[RocketCore.scala 743:54]
  assign _T_1675 = io_fpu_dec_ren1 & _T_1666; // @[RocketCore.scala 983:27]
  assign _T_1677 = io_fpu_dec_ren2 & _T_1668; // @[RocketCore.scala 983:27]
  assign _T_1682 = _T_1675 | _T_1677; // @[RocketCore.scala 983:50]
  assign _T_1678 = id_raddr3 == wb_waddr; // @[RocketCore.scala 742:76]
  assign _T_1679 = io_fpu_dec_ren3 & _T_1678; // @[RocketCore.scala 983:27]
  assign _T_1683 = _T_1682 | _T_1679; // @[RocketCore.scala 983:50]
  assign _T_1681 = io_fpu_dec_wen & _T_1670; // @[RocketCore.scala 983:27]
  assign _T_1684 = _T_1683 | _T_1681; // @[RocketCore.scala 983:50]
  assign fp_data_hazard_wb = wb_ctrl_wfd & _T_1684; // @[RocketCore.scala 742:39]
  assign _T_1686 = _T_1685 | fp_data_hazard_wb; // @[RocketCore.scala 743:71]
  assign id_wb_hazard = wb_reg_valid & _T_1686; // @[RocketCore.scala 743:35]
  assign _T_1734 = _T_1733 | id_wb_hazard; // @[RocketCore.scala 764:35]
  assign _T_1576 = {_T_1574[31:1], 1'h0}; // @[RocketCore.scala 1001:40]
  assign _T_1582 = _T_1576 >> id_raddr1; // @[RocketCore.scala 997:35]
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data; // @[RocketCore.scala 638:44]
  assign dmem_resp_replay = dmem_resp_valid & io_dmem_resp_bits_replay; // @[RocketCore.scala 639:42]
  assign dmem_resp_xpu = ~io_dmem_resp_bits_tag[0]; // @[RocketCore.scala 635:23]
  assign _T_1511 = dmem_resp_replay & dmem_resp_xpu; // @[RocketCore.scala 654:26]
  assign _T_1510 = div_io_resp_ready & div_io_resp_valid; // @[Decoupled.scala 40:37]
  assign ll_wen = _T_1511 | _T_1510; // @[RocketCore.scala 654:44]
  assign dmem_resp_waddr = io_dmem_resp_bits_tag[5:1]; // @[RocketCore.scala 637:46]
  assign ll_waddr = _T_1511 ? dmem_resp_waddr : div_io_resp_bits_tag; // @[RocketCore.scala 654:44]
  assign _T_1584 = ll_waddr == id_raddr1; // @[RocketCore.scala 718:70]
  assign _T_1585 = ll_wen & _T_1584; // @[RocketCore.scala 718:58]
  assign _T_1587 = _T_1582[0] & ~_T_1585; // @[RocketCore.scala 721:77]
  assign _T_1588 = _T_1569 & _T_1587; // @[RocketCore.scala 983:27]
  assign _T_1589 = _T_1576 >> id_raddr2; // @[RocketCore.scala 997:35]
  assign _T_1591 = ll_waddr == id_raddr2; // @[RocketCore.scala 718:70]
  assign _T_1592 = ll_wen & _T_1591; // @[RocketCore.scala 718:58]
  assign _T_1594 = _T_1589[0] & ~_T_1592; // @[RocketCore.scala 721:77]
  assign _T_1595 = _T_1571 & _T_1594; // @[RocketCore.scala 983:27]
  assign _T_1603 = _T_1588 | _T_1595; // @[RocketCore.scala 983:50]
  assign _T_1596 = _T_1576 >> id_waddr; // @[RocketCore.scala 997:35]
  assign _T_1598 = ll_waddr == id_waddr; // @[RocketCore.scala 718:70]
  assign _T_1599 = ll_wen & _T_1598; // @[RocketCore.scala 718:58]
  assign _T_1601 = _T_1596[0] & ~_T_1599; // @[RocketCore.scala 721:77]
  assign _T_1602 = _T_1573 & _T_1601; // @[RocketCore.scala 983:27]
  assign id_sboard_hazard = _T_1603 | _T_1602; // @[RocketCore.scala 983:50]
  assign _T_1735 = _T_1734 | id_sboard_hazard; // @[RocketCore.scala 764:51]
  assign _T_1736 = ex_reg_valid | mem_reg_valid; // @[RocketCore.scala 765:40]
  assign _T_1737 = _T_1736 | wb_reg_valid; // @[RocketCore.scala 765:57]
  assign _T_1738 = csr_io_singleStep & _T_1737; // @[RocketCore.scala 765:23]
  assign _T_1739 = _T_1735 | _T_1738; // @[RocketCore.scala 764:71]
  assign _T_1740 = id_csr_en & csr_io_decode_0_fp_csr; // @[RocketCore.scala 766:15]
  assign _T_1742 = _T_1740 & ~io_fpu_fcsr_rdy; // @[RocketCore.scala 766:42]
  assign _T_1743 = _T_1739 | _T_1742; // @[RocketCore.scala 765:74]
  assign _T_1706 = _T_1687 >> id_raddr1; // @[RocketCore.scala 997:35]
  assign _T_1708 = io_fpu_dec_ren1 & _T_1706[0]; // @[RocketCore.scala 983:27]
  assign _T_1709 = _T_1687 >> id_raddr2; // @[RocketCore.scala 997:35]
  assign _T_1711 = io_fpu_dec_ren2 & _T_1709[0]; // @[RocketCore.scala 983:27]
  assign _T_1718 = _T_1708 | _T_1711; // @[RocketCore.scala 983:50]
  assign _T_1712 = _T_1687 >> id_raddr3; // @[RocketCore.scala 997:35]
  assign _T_1714 = io_fpu_dec_ren3 & _T_1712[0]; // @[RocketCore.scala 983:27]
  assign _T_1719 = _T_1718 | _T_1714; // @[RocketCore.scala 983:50]
  assign _T_1715 = _T_1687 >> id_waddr; // @[RocketCore.scala 997:35]
  assign _T_1717 = io_fpu_dec_wen & _T_1715[0]; // @[RocketCore.scala 983:27]
  assign id_stall_fpu = _T_1719 | _T_1717; // @[RocketCore.scala 983:50]
  assign _T_1744 = id_ctrl_fp & id_stall_fpu; // @[RocketCore.scala 767:16]
  assign _T_1745 = _T_1743 | _T_1744; // @[RocketCore.scala 766:62]
  assign dcache_blocked = blocked & ~io_dmem_perf_grant; // @[RocketCore.scala 758:13]
  assign _T_1746 = id_ctrl_mem & dcache_blocked; // @[RocketCore.scala 768:17]
  assign _T_1747 = _T_1745 | _T_1746; // @[RocketCore.scala 767:32]
  assign wb_wxd = wb_reg_valid & wb_ctrl_wxd; // @[RocketCore.scala 627:29]
  assign _T_1751 = div_io_resp_valid & ~wb_wxd; // @[RocketCore.scala 770:62]
  assign _T_1752 = div_io_req_ready | _T_1751; // @[RocketCore.scala 770:40]
  assign _T_1754 = ~_T_1752 | div_io_req_valid; // @[RocketCore.scala 770:75]
  assign _T_1755 = id_ctrl_div & _T_1754; // @[RocketCore.scala 770:17]
  assign _T_1756 = _T_1747 | _T_1755; // @[RocketCore.scala 769:34]
  assign _T_1759 = _T_1756 | id_do_fence; // @[RocketCore.scala 771:15]
  assign _T_1760 = _T_1759 | csr_io_csr_stall; // @[RocketCore.scala 772:17]
  assign ctrl_stalld = _T_1760 | id_reg_pause; // @[RocketCore.scala 773:22]
  assign _T_1765 = _T_1764 | ctrl_stalld; // @[RocketCore.scala 776:89]
  assign ctrl_killd = _T_1765 | csr_io_interrupt; // @[RocketCore.scala 776:104]
  assign _T_1102 = ~take_pc_mem_wb & ibuf_io_inst_0_valid; // @[RocketCore.scala 416:29]
  assign _T_1112 = id_fence_succ == 4'h0; // @[RocketCore.scala 426:42]
  assign _T_1113 = id_ctrl_fence & _T_1112; // @[RocketCore.scala 426:25]
  assign _GEN_1 = _T_1113 | id_reg_pause; // @[RocketCore.scala 426:49]
  assign _GEN_2 = id_fence_next | _GEN_0; // @[RocketCore.scala 427:26]
  assign _T_1114 = {ibuf_io_inst_0_bits_xcpt1_pf_inst,ibuf_io_inst_0_bits_xcpt1_ae_inst}; // @[RocketCore.scala 433:22]
  assign _T_1115 = |_T_1114; // @[RocketCore.scala 433:29]
  assign _GEN_5 = _T_1115 | ibuf_io_inst_0_bits_rvc; // @[RocketCore.scala 433:34]
  assign _T_1116 = {ibuf_io_inst_0_bits_xcpt0_pf_inst,ibuf_io_inst_0_bits_xcpt0_ae_inst}; // @[RocketCore.scala 438:40]
  assign _T_1117 = |_T_1116; // @[RocketCore.scala 438:47]
  assign _T_1118 = bpu_io_xcpt_if | _T_1117; // @[RocketCore.scala 438:28]
  assign _GEN_9 = id_xcpt | id_ctrl_alu_dw; // @[RocketCore.scala 428:20]
  assign _T_1119 = id_ctrl_fence_i | id_csr_flush; // @[RocketCore.scala 443:42]
  assign _T_1122 = id_ctrl_mem_cmd == 5'h5; // @[package.scala 15:47]
  assign _T_1123 = _T_902 | _T_1122; // @[package.scala 64:59]
  assign _T_1126 = {_T_1570,_T_1568}; // @[Cat.scala 29:58]
  assign _T_1127 = id_bypass_src_0_0 | id_bypass_src_0_1; // @[RocketCore.scala 456:48]
  assign _T_1128 = _T_1127 | id_bypass_src_0_2; // @[RocketCore.scala 456:48]
  assign do_bypass = _T_1128 | id_bypass_src_0_3; // @[RocketCore.scala 456:48]
  assign _T_1132 = id_ctrl_rxs1 & ~do_bypass; // @[RocketCore.scala 460:23]
  assign _T_1513 = wb_reg_valid & ~replay_wb_common; // @[RocketCore.scala 662:31]
  assign wb_valid = _T_1513 & ~wb_xcpt; // @[RocketCore.scala 662:45]
  assign wb_wen = wb_valid & wb_ctrl_wxd; // @[RocketCore.scala 663:25]
  assign rf_wen = wb_wen | ll_wen; // @[RocketCore.scala 664:23]
  assign rf_waddr = ll_wen ? ll_waddr : wb_waddr; // @[RocketCore.scala 665:21]
  assign _T_1521 = rf_waddr != 5'h0; // @[RocketCore.scala 1026:16]
  assign _T_1525 = rf_waddr == id_raddr1; // @[RocketCore.scala 1029:20]
  assign _T_1515 = dmem_resp_valid & dmem_resp_xpu; // @[RocketCore.scala 666:38]
  assign ll_wdata = div_io_resp_bits_data;
  assign _T_1517 = wb_ctrl_csr != 3'h0; // @[RocketCore.scala 668:34]
  assign _T_1519 = _T_1517 ? csr_io_rw_rdata : wb_reg_wdata; // @[RocketCore.scala 668:21]
  assign _T_1520 = ll_wen ? ll_wdata : _T_1519; // @[RocketCore.scala 667:21]
  assign rf_wdata = _T_1515 ? io_dmem_resp_bits_data : _T_1520; // @[RocketCore.scala 666:21]
  assign _GEN_226 = _T_1525 ? rf_wdata : _T_821; // @[RocketCore.scala 1029:31]
  assign _GEN_233 = _T_1521 ? _GEN_226 : _T_821; // @[RocketCore.scala 1026:29]
  assign id_rs_0 = rf_wen ? _GEN_233 : _T_821; // @[RocketCore.scala 671:17]
  assign _T_1135 = id_bypass_src_1_0 | id_bypass_src_1_1; // @[RocketCore.scala 456:48]
  assign _T_1136 = _T_1135 | id_bypass_src_1_2; // @[RocketCore.scala 456:48]
  assign do_bypass_1 = _T_1136 | id_bypass_src_1_3; // @[RocketCore.scala 456:48]
  assign _T_1140 = id_ctrl_rxs2 & ~do_bypass_1; // @[RocketCore.scala 460:23]
  assign _T_1526 = rf_waddr == id_raddr2; // @[RocketCore.scala 1029:20]
  assign _GEN_227 = _T_1526 ? rf_wdata : _T_827; // @[RocketCore.scala 1029:31]
  assign _GEN_234 = _T_1521 ? _GEN_227 : _T_827; // @[RocketCore.scala 1026:29]
  assign id_rs_1 = rf_wen ? _GEN_234 : _T_827; // @[RocketCore.scala 671:17]
  assign inst = ibuf_io_inst_0_bits_rvc ? {{16'd0}, ibuf_io_inst_0_bits_raw[15:0]} : ibuf_io_inst_0_bits_raw; // @[RocketCore.scala 466:21]
  assign _T_1664 = mem_reg_valid & data_hazard_mem; // @[RocketCore.scala 738:32]
  assign id_load_use = _T_1664 & mem_ctrl_mem; // @[RocketCore.scala 738:51]
  assign _T_1147 = ~ctrl_killd | csr_io_interrupt; // @[RocketCore.scala 472:21]
  assign _T_1148 = _T_1147 | ibuf_io_inst_0_bits_replay; // @[RocketCore.scala 472:41]
  assign _T_1152 = ex_ctrl_mem & ~io_dmem_req_ready; // @[RocketCore.scala 484:42]
  assign _T_1154 = ex_ctrl_div & ~div_io_req_ready; // @[RocketCore.scala 485:42]
  assign replay_ex_structural = _T_1152 | _T_1154; // @[RocketCore.scala 484:64]
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use; // @[RocketCore.scala 486:43]
  assign _T_1155 = replay_ex_structural | replay_ex_load_use; // @[RocketCore.scala 487:75]
  assign _T_1156 = ex_reg_valid & _T_1155; // @[RocketCore.scala 487:50]
  assign replay_ex = ex_reg_replay | _T_1156; // @[RocketCore.scala 487:33]
  assign _T_1157 = take_pc_mem_wb | replay_ex; // @[RocketCore.scala 488:35]
  assign ctrl_killx = _T_1157 | ~ex_reg_valid; // @[RocketCore.scala 488:48]
  assign _T_1159 = ex_ctrl_mem_cmd == 5'h7; // @[RocketCore.scala 490:40]
  assign _T_1160 = ex_reg_mem_size < 2'h2; // @[RocketCore.scala 490:69]
  assign ex_slow_bypass = _T_1159 | _T_1160; // @[RocketCore.scala 490:50]
  assign _T_1162 = ex_ctrl_mem_cmd == 5'h14; // @[RocketCore.scala 491:67]
  assign ex_sfence = ex_ctrl_mem & _T_1162; // @[RocketCore.scala 491:48]
  assign ex_xcpt = ex_reg_xcpt_interrupt | ex_reg_xcpt; // @[RocketCore.scala 494:28]
  assign _T_1173 = mem_reg_valid | mem_reg_replay; // @[RocketCore.scala 500:36]
  assign mem_pc_valid = _T_1173 | mem_reg_xcpt_interrupt; // @[RocketCore.scala 500:54]
  assign _T_1326 = ~csr_io_status_isa[2] & mem_npc[1]; // @[RocketCore.scala 509:56]
  assign mem_npc_misaligned = _T_1326 & ~mem_reg_sfence; // @[RocketCore.scala 509:70]
  assign _T_1329 = mem_ctrl_jalr ^ mem_npc_misaligned; // @[RocketCore.scala 510:59]
  assign _T_1330 = ~mem_reg_xcpt & _T_1329; // @[RocketCore.scala 510:41]
  assign mem_int_wdata = _T_1330 ? $signed({{24{mem_br_target[39]}},mem_br_target}) : $signed(mem_reg_wdata); // @[RocketCore.scala 510:119]
  assign _T_1333 = mem_ctrl_branch | mem_ctrl_jalr; // @[RocketCore.scala 511:33]
  assign mem_cfi = _T_1333 | mem_ctrl_jal; // @[RocketCore.scala 511:50]
  assign _T_1335 = _T_1175 | mem_ctrl_jalr; // @[RocketCore.scala 512:57]
  assign mem_cfi_taken = _T_1335 | mem_ctrl_jal; // @[RocketCore.scala 512:74]
  assign _T_1347 = mem_reg_valid & mem_reg_flush_pipe; // @[RocketCore.scala 524:23]
  assign _T_1348 = ex_ctrl_mem_cmd == 5'h0; // @[Consts.scala 82:31]
  assign _T_1349 = ex_ctrl_mem_cmd == 5'h6; // @[Consts.scala 82:48]
  assign _T_1350 = _T_1348 | _T_1349; // @[Consts.scala 82:41]
  assign _T_1352 = _T_1350 | _T_1159; // @[Consts.scala 82:58]
  assign _T_1353 = ex_ctrl_mem_cmd == 5'h4; // @[package.scala 15:47]
  assign _T_1354 = ex_ctrl_mem_cmd == 5'h9; // @[package.scala 15:47]
  assign _T_1355 = ex_ctrl_mem_cmd == 5'ha; // @[package.scala 15:47]
  assign _T_1356 = ex_ctrl_mem_cmd == 5'hb; // @[package.scala 15:47]
  assign _T_1357 = _T_1353 | _T_1354; // @[package.scala 64:59]
  assign _T_1358 = _T_1357 | _T_1355; // @[package.scala 64:59]
  assign _T_1359 = _T_1358 | _T_1356; // @[package.scala 64:59]
  assign _T_1360 = ex_ctrl_mem_cmd == 5'h8; // @[package.scala 15:47]
  assign _T_1361 = ex_ctrl_mem_cmd == 5'hc; // @[package.scala 15:47]
  assign _T_1362 = ex_ctrl_mem_cmd == 5'hd; // @[package.scala 15:47]
  assign _T_1363 = ex_ctrl_mem_cmd == 5'he; // @[package.scala 15:47]
  assign _T_1364 = ex_ctrl_mem_cmd == 5'hf; // @[package.scala 15:47]
  assign _T_1365 = _T_1360 | _T_1361; // @[package.scala 64:59]
  assign _T_1366 = _T_1365 | _T_1362; // @[package.scala 64:59]
  assign _T_1367 = _T_1366 | _T_1363; // @[package.scala 64:59]
  assign _T_1368 = _T_1367 | _T_1364; // @[package.scala 64:59]
  assign _T_1369 = _T_1359 | _T_1368; // @[Consts.scala 80:44]
  assign _T_1370 = _T_1352 | _T_1369; // @[Consts.scala 82:75]
  assign _T_1371 = ex_ctrl_mem & _T_1370; // @[RocketCore.scala 531:33]
  assign _T_1372 = ex_ctrl_mem_cmd == 5'h1; // @[Consts.scala 83:32]
  assign _T_1373 = ex_ctrl_mem_cmd == 5'h11; // @[Consts.scala 83:49]
  assign _T_1374 = _T_1372 | _T_1373; // @[Consts.scala 83:42]
  assign _T_1376 = _T_1374 | _T_1159; // @[Consts.scala 83:59]
  assign _T_1394 = _T_1376 | _T_1369; // @[Consts.scala 83:76]
  assign _T_1395 = ex_ctrl_mem & _T_1394; // @[RocketCore.scala 532:34]
  assign _T_1396 = alu_io_out; // @[RocketCore.scala 544:25]
  assign _T_1398 = ex_ctrl_mem | ex_sfence; // @[RocketCore.scala 547:56]
  assign _T_1399 = ex_ctrl_rxs2 & _T_1398; // @[RocketCore.scala 547:24]
  assign _T_1401 = ex_reg_mem_size == 2'h0; // @[AMOALU.scala 26:19]
  assign _T_1405 = {ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[7:0]}; // @[Cat.scala 29:58]
  assign _T_1406 = ex_reg_mem_size == 2'h1; // @[AMOALU.scala 26:19]
  assign _T_1409 = {ex_rs_1[15:0],ex_rs_1[15:0],ex_rs_1[15:0],ex_rs_1[15:0]}; // @[Cat.scala 29:58]
  assign _T_1410 = ex_reg_mem_size == 2'h2; // @[AMOALU.scala 26:19]
  assign _T_1412 = {ex_rs_1[31:0],ex_rs_1[31:0]}; // @[Cat.scala 29:58]
  assign _T_1416 = ex_ctrl_jalr & csr_io_status_debug; // @[RocketCore.scala 551:24]
  assign _GEN_77 = _T_1416 | ex_ctrl_fence_i; // @[RocketCore.scala 551:48]
  assign _GEN_78 = _T_1416 | ex_reg_flush_pipe; // @[RocketCore.scala 551:48]
  assign _T_1417 = mem_reg_load & bpu_io_xcpt_ld; // @[RocketCore.scala 558:38]
  assign _T_1418 = mem_reg_store & bpu_io_xcpt_st; // @[RocketCore.scala 558:75]
  assign mem_breakpoint = _T_1417 | _T_1418; // @[RocketCore.scala 558:57]
  assign _T_1419 = mem_reg_load & bpu_io_debug_ld; // @[RocketCore.scala 559:44]
  assign _T_1420 = mem_reg_store & bpu_io_debug_st; // @[RocketCore.scala 559:82]
  assign mem_debug_breakpoint = _T_1419 | _T_1420; // @[RocketCore.scala 559:64]
  assign mem_ldst_xcpt = mem_debug_breakpoint | mem_breakpoint; // @[RocketCore.scala 974:26]
  assign mem_ldst_cause = mem_debug_breakpoint ? 4'he : 4'h3; // @[Mux.scala 47:69]
  assign _T_1421 = mem_reg_xcpt_interrupt | mem_reg_xcpt; // @[RocketCore.scala 565:29]
  assign _T_1422 = mem_reg_valid & mem_npc_misaligned; // @[RocketCore.scala 566:20]
  assign _T_1423 = mem_reg_valid & mem_ldst_xcpt; // @[RocketCore.scala 567:20]
  assign _T_1424 = _T_1421 | _T_1422; // @[RocketCore.scala 974:26]
  assign mem_xcpt = _T_1424 | _T_1423; // @[RocketCore.scala 974:26]
  assign _T_1425 = _T_1422 ? 4'h0 : mem_ldst_cause; // @[Mux.scala 47:69]
  assign dcache_kill_mem = _T_998 & io_dmem_replay_next; // @[RocketCore.scala 576:55]
  assign _T_1439 = mem_reg_valid & mem_ctrl_fp; // @[RocketCore.scala 577:36]
  assign fpu_kill_mem = _T_1439 & io_fpu_nack_mem; // @[RocketCore.scala 577:51]
  assign _T_1440 = dcache_kill_mem | mem_reg_replay; // @[RocketCore.scala 578:37]
  assign replay_mem = _T_1440 | fpu_kill_mem; // @[RocketCore.scala 578:55]
  assign _T_1441 = dcache_kill_mem | take_pc_wb; // @[RocketCore.scala 579:38]
  assign _T_1442 = _T_1441 | mem_reg_xcpt; // @[RocketCore.scala 579:52]
  assign killm_common = _T_1442 | ~mem_reg_valid; // @[RocketCore.scala 579:68]
  assign _T_1447 = killm_common | mem_xcpt; // @[RocketCore.scala 581:33]
  assign ctrl_killm = _T_1447 | fpu_kill_mem; // @[RocketCore.scala 581:45]
  assign _T_1456 = ~mem_reg_xcpt & mem_ctrl_fp; // @[RocketCore.scala 592:25]
  assign _T_1457 = _T_1456 & mem_ctrl_wxd; // @[RocketCore.scala 592:40]
  assign _T_1482 = _T_1474 ? 3'h7 : 3'h5; // @[Mux.scala 47:69]
  assign _T_1483 = _T_1472 ? 4'hd : {{1'd0}, _T_1482}; // @[Mux.scala 47:69]
  assign _T_1484 = _T_1470 ? 4'hf : _T_1483; // @[Mux.scala 47:69]
  assign _T_1485 = _T_1468 ? 4'h4 : _T_1484; // @[Mux.scala 47:69]
  assign _T_1486 = _T_1466 ? 4'h6 : _T_1485; // @[Mux.scala 47:69]
  assign wb_cause = wb_reg_xcpt ? wb_reg_cause : {{60'd0}, _T_1486}; // @[Mux.scala 47:69]
  assign _T_1487 = wb_cause == 64'h6; // @[RocketCore.scala 978:38]
  assign _T_1489 = wb_cause == 64'h4; // @[RocketCore.scala 978:38]
  assign _T_1491 = wb_cause == 64'h7; // @[RocketCore.scala 978:38]
  assign _T_1493 = wb_cause == 64'h5; // @[RocketCore.scala 978:38]
  assign _T_1495 = wb_cause == 64'hf; // @[RocketCore.scala 978:38]
  assign _T_1497 = wb_cause == 64'hd; // @[RocketCore.scala 978:38]
  assign _T_1529 = &wb_reg_raw_inst[1:0]; // @[RocketCore.scala 679:73]
  assign _T_1531 = _T_1529 ? wb_reg_inst[31:16] : 16'h0; // @[RocketCore.scala 679:50]
  assign _T_1535 = wb_cause == 64'h2; // @[package.scala 15:47]
  assign _T_1536 = wb_cause == 64'h3; // @[package.scala 15:47]
  assign _T_1541 = wb_cause == 64'h1; // @[package.scala 15:47]
  assign _T_1544 = wb_cause == 64'hc; // @[package.scala 15:47]
  assign _T_1545 = _T_1535 | _T_1536; // @[package.scala 64:59]
  assign _T_1546 = _T_1545 | _T_1489; // @[package.scala 64:59]
  assign _T_1547 = _T_1546 | _T_1487; // @[package.scala 64:59]
  assign _T_1548 = _T_1547 | _T_1493; // @[package.scala 64:59]
  assign _T_1549 = _T_1548 | _T_1491; // @[package.scala 64:59]
  assign _T_1550 = _T_1549 | _T_1541; // @[package.scala 64:59]
  assign _T_1551 = _T_1550 | _T_1497; // @[package.scala 64:59]
  assign _T_1552 = _T_1551 | _T_1495; // @[package.scala 64:59]
  assign _T_1553 = _T_1552 | _T_1544; // @[package.scala 64:59]
  assign tval_valid = wb_xcpt & _T_1553; // @[RocketCore.scala 688:28]
  assign a_1 = wb_reg_wdata[63:39]; // @[RocketCore.scala 988:23]
  assign _T_1555 = $signed(a_1) == 25'sh0; // @[RocketCore.scala 989:21]
  assign _T_1556 = $signed(a_1) == -25'sh1; // @[RocketCore.scala 989:34]
  assign _T_1557 = _T_1555 | _T_1556; // @[RocketCore.scala 989:29]
  assign msb_1 = _T_1557 ? wb_reg_wdata[39] : ~wb_reg_wdata[38]; // @[RocketCore.scala 989:18]
  assign _T_1562 = {msb_1,wb_reg_wdata[38:0]}; // @[Cat.scala 29:58]
  assign _T_1565 = wb_reg_valid ? 3'h0 : 3'h4; // @[CSR.scala 131:15]
  assign _T_1577 = 32'h1 << ll_waddr; // @[RocketCore.scala 1004:62]
  assign _T_1578 = ll_wen ? _T_1577 : 32'h0; // @[RocketCore.scala 1004:49]
  assign _T_1580 = _T_1576 & ~_T_1578; // @[RocketCore.scala 996:62]
  assign _T_1604 = wb_set_sboard & wb_wen; // @[RocketCore.scala 722:28]
  assign _T_1605 = 32'h1 << wb_waddr; // @[RocketCore.scala 1004:62]
  assign _T_1606 = _T_1604 ? _T_1605 : 32'h0; // @[RocketCore.scala 1004:49]
  assign _T_1607 = _T_1580 | _T_1606; // @[RocketCore.scala 995:60]
  assign _T_1608 = ll_wen | _T_1604; // @[RocketCore.scala 1007:17]
  assign _T_1688 = wb_dcache_miss & wb_ctrl_wfd; // @[RocketCore.scala 747:35]
  assign _T_1689 = _T_1688 | io_fpu_sboard_set; // @[RocketCore.scala 747:50]
  assign _T_1690 = _T_1689 & wb_valid; // @[RocketCore.scala 747:72]
  assign _T_1692 = _T_1690 ? _T_1605 : 32'h0; // @[RocketCore.scala 1004:49]
  assign _T_1693 = _T_1687 | _T_1692; // @[RocketCore.scala 995:60]
  assign _T_1695 = dmem_resp_replay & io_dmem_resp_bits_tag[0]; // @[RocketCore.scala 748:38]
  assign _T_1696 = 32'h1 << dmem_resp_waddr; // @[RocketCore.scala 1004:62]
  assign _T_1697 = _T_1695 ? _T_1696 : 32'h0; // @[RocketCore.scala 1004:49]
  assign _T_1699 = _T_1693 & ~_T_1697; // @[RocketCore.scala 996:62]
  assign _T_1700 = _T_1690 | _T_1695; // @[RocketCore.scala 1007:17]
  assign _T_1701 = 32'h1 << io_fpu_sboard_clra; // @[RocketCore.scala 1004:62]
  assign _T_1702 = io_fpu_sboard_clr ? _T_1701 : 32'h0; // @[RocketCore.scala 1004:49]
  assign _T_1704 = _T_1699 & ~_T_1702; // @[RocketCore.scala 996:62]
  assign _T_1705 = _T_1700 | io_fpu_sboard_clr; // @[RocketCore.scala 1007:17]
  assign _T_1723 = ~io_dmem_req_ready & ~io_dmem_perf_grant; // @[RocketCore.scala 757:60]
  assign _T_1724 = blocked | io_dmem_req_valid; // @[RocketCore.scala 757:95]
  assign _T_1725 = _T_1724 | io_dmem_s2_nack; // @[RocketCore.scala 757:116]
  assign _T_1768 = wb_xcpt | csr_io_eret; // @[RocketCore.scala 781:17]
  assign _T_1769 = replay_wb_common ? wb_reg_pc : mem_npc; // @[RocketCore.scala 782:8]
  assign _T_1771 = wb_reg_valid & wb_ctrl_fence_i; // @[RocketCore.scala 784:40]
  assign _T_1774 = ex_pc_valid | mem_pc_valid; // @[RocketCore.scala 786:43]
  assign _T_1782 = mem_reg_valid & ~take_pc_wb; // @[RocketCore.scala 798:45]
  assign _T_1783 = _T_1782 & mem_wrong_npc; // @[RocketCore.scala 798:60]
  assign _T_1785 = ~mem_cfi | mem_cfi_taken; // @[RocketCore.scala 798:90]
  assign _T_1787 = mem_ctrl_jal | mem_ctrl_jalr; // @[RocketCore.scala 801:23]
  assign _T_1789 = _T_1787 & mem_waddr[0]; // @[RocketCore.scala 801:41]
  assign _T_1792 = mem_reg_inst[19:15] & 5'h1b; // @[RocketCore.scala 802:62]
  assign _T_1793 = 5'h1 == _T_1792; // @[RocketCore.scala 802:62]
  assign _T_1794 = mem_ctrl_jalr & _T_1793; // @[RocketCore.scala 802:23]
  assign _T_1797 = _T_1794 ? 2'h3 : {{1'd0}, _T_1787}; // @[RocketCore.scala 802:8]
  assign _T_1799 = mem_reg_rvc ? 2'h0 : 2'h2; // @[RocketCore.scala 806:74]
  assign _GEN_250 = {{38'd0}, _T_1799}; // @[RocketCore.scala 806:69]
  assign _T_1801 = mem_reg_pc + _GEN_250; // @[RocketCore.scala 806:69]
  assign _T_1803 = ~io_imem_btb_update_bits_br_pc | 39'h3; // @[RocketCore.scala 807:66]
  assign ex_dcache_tag = {ex_waddr,ex_ctrl_fp}; // @[Cat.scala 29:58]
  assign a_2 = _T_1085[63:39]; // @[RocketCore.scala 988:23]
  assign _T_1815 = $signed(a_2) == 25'sh0; // @[RocketCore.scala 989:21]
  assign _T_1816 = $signed(a_2) == -25'sh1; // @[RocketCore.scala 989:34]
  assign _T_1817 = _T_1815 | _T_1816; // @[RocketCore.scala 989:29]
  assign msb_2 = _T_1817 ? alu_io_adder_out[39] : ~alu_io_adder_out[38]; // @[RocketCore.scala 989:18]
  assign _T_1824 = killm_common | mem_ldst_xcpt; // @[RocketCore.scala 839:35]
  assign _T_1845 = csr_io_time[4:0] == 5'h0; // @[RocketCore.scala 852:62]
  assign _T_1846 = _T_1845 | io_dmem_perf_release; // @[RocketCore.scala 852:68]
  assign unpause = _T_1846 | take_pc_mem_wb; // @[RocketCore.scala 852:92]
  assign _T_1849 = ibuf_io_inst_0_ready & ibuf_io_inst_0_valid; // @[RocketCore.scala 871:33]
  assign coreMonitorBundle_valid = csr_io_trace_0_valid & ~csr_io_trace_0_exception; // @[RocketCore.scala 888:52]
  assign _T_1858 = csr_io_trace_0_iaddr; // @[RocketCore.scala 889:48]
  assign _T_1861 = _T_1858[39] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign coreMonitorBundle_pc = {_T_1861,_T_1858}; // @[Cat.scala 29:58]
  assign coreMonitorBundle_wrenx = wb_wen & ~wb_set_sboard; // @[RocketCore.scala 890:37]
  assign _T_1871 = wb_ctrl_wxd | wb_ctrl_wfd; // @[RocketCore.scala 933:26]
  assign _T_1872 = _T_1871 ? wb_waddr : 5'h0; // @[RocketCore.scala 933:13]
  assign _T_1873 = coreMonitorBundle_wrenx ? rf_wdata : 64'h0; // @[RocketCore.scala 934:13]
  assign _T_1874 = wb_ctrl_rxs1 | wb_ctrl_rfs1; // @[RocketCore.scala 936:27]
  assign _T_1875 = _T_1874 ? wb_reg_inst[19:15] : 5'h0; // @[RocketCore.scala 936:13]
  assign _T_1877 = _T_1874 ? coreMonitorBundle_rd0val : 64'h0; // @[RocketCore.scala 937:13]
  assign _T_1878 = wb_ctrl_rxs2 | wb_ctrl_rfs2; // @[RocketCore.scala 938:27]
  assign _T_1879 = _T_1878 ? wb_reg_inst[24:20] : 5'h0; // @[RocketCore.scala 938:13]
  assign _T_1881 = _T_1878 ? coreMonitorBundle_rd1val : 64'h0; // @[RocketCore.scala 939:13]
  assign coreMonitorBundle_inst = csr_io_trace_0_insn; // @[RocketCore.scala 882:31 RocketCore.scala 898:26]
  assign io_imem_might_request = imem_might_request_reg; // @[RocketCore.scala 785:25]
  assign io_imem_req_valid = take_pc_wb | take_pc_mem; // @[RocketCore.scala 778:21]
  assign io_imem_req_bits_pc = _T_1768 ? csr_io_evec : _T_1769; // @[RocketCore.scala 780:23]
  assign io_imem_req_bits_speculative = ~take_pc_wb; // @[RocketCore.scala 779:32]
  assign io_imem_sfence_valid = wb_reg_valid & wb_reg_sfence; // @[RocketCore.scala 789:24]
  assign io_imem_sfence_bits_rs1 = wb_reg_mem_size[0]; // @[RocketCore.scala 790:27]
  assign io_imem_sfence_bits_rs2 = wb_reg_mem_size[1]; // @[RocketCore.scala 791:27]
  assign io_imem_sfence_bits_addr = wb_reg_wdata[38:0]; // @[RocketCore.scala 792:28]
  assign io_imem_resp_ready = ibuf_io_imem_ready; // @[RocketCore.scala 252:16]
  assign io_imem_btb_update_valid = _T_1783 & _T_1785; // @[RocketCore.scala 798:28]
  assign io_imem_btb_update_bits_prediction_entry = mem_reg_btb_resp_entry; // @[RocketCore.scala 808:38]
  assign io_imem_btb_update_bits_pc = ~_T_1803; // @[RocketCore.scala 807:30]
  assign io_imem_btb_update_bits_isValid = _T_1333 | mem_ctrl_jal; // @[RocketCore.scala 799:35]
  assign io_imem_btb_update_bits_br_pc = _T_1801[38:0]; // @[RocketCore.scala 806:33]
  assign io_imem_btb_update_bits_cfiType = _T_1789 ? 2'h2 : _T_1797; // @[RocketCore.scala 800:35]
  assign io_imem_bht_update_valid = mem_reg_valid & ~take_pc_wb; // @[RocketCore.scala 810:28]
  assign io_imem_bht_update_bits_prediction_history = mem_reg_btb_resp_bht_history; // @[RocketCore.scala 815:38]
  assign io_imem_bht_update_bits_pc = io_imem_btb_update_bits_pc; // @[RocketCore.scala 811:30]
  assign io_imem_bht_update_bits_branch = mem_ctrl_branch; // @[RocketCore.scala 814:34]
  assign io_imem_bht_update_bits_taken = mem_br_taken; // @[RocketCore.scala 812:33]
  assign io_imem_bht_update_bits_mispredict = ex_pc_valid ? _T_1319 : _T_1322; // @[RocketCore.scala 813:38]
  assign io_imem_flush_icache = _T_1771 & ~io_dmem_s2_nack; // @[RocketCore.scala 784:24]
  assign io_dmem_req_valid = ex_reg_valid & ex_ctrl_mem; // @[RocketCore.scala 828:25]
  assign io_dmem_req_bits_addr = {msb_2,alu_io_adder_out[38:0]}; // @[RocketCore.scala 836:25]
  assign io_dmem_req_bits_tag = {{1'd0}, ex_dcache_tag}; // @[RocketCore.scala 831:25]
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd; // @[RocketCore.scala 832:25]
  assign io_dmem_req_bits_size = ex_reg_mem_size; // @[RocketCore.scala 833:25]
  assign io_dmem_req_bits_signed = ~ex_reg_inst[14]; // @[RocketCore.scala 834:27]
  assign io_dmem_s1_kill = _T_1824 | fpu_kill_mem; // @[RocketCore.scala 839:19]
  assign io_dmem_s1_data_data = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2; // @[RocketCore.scala 838:24]
  assign io_ptw_ptbr_mode = csr_io_ptbr_mode; // @[RocketCore.scala 693:15]
  assign io_ptw_ptbr_ppn = csr_io_ptbr_ppn; // @[RocketCore.scala 693:15]
  assign io_ptw_sfence_valid = io_imem_sfence_valid; // @[RocketCore.scala 794:17]
  assign io_ptw_sfence_bits_rs1 = io_imem_sfence_bits_rs1; // @[RocketCore.scala 794:17]
  assign io_ptw_status_debug = csr_io_status_debug; // @[RocketCore.scala 695:17]
  assign io_ptw_status_dprv = csr_io_status_dprv; // @[RocketCore.scala 695:17]
  assign io_ptw_status_prv = csr_io_status_prv; // @[RocketCore.scala 695:17]
  assign io_ptw_status_mxr = csr_io_status_mxr; // @[RocketCore.scala 695:17]
  assign io_ptw_status_sum = csr_io_status_sum; // @[RocketCore.scala 695:17]
  assign io_ptw_pmp_0_cfg_l = csr_io_pmp_0_cfg_l; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_0_cfg_a = csr_io_pmp_0_cfg_a; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_0_cfg_x = csr_io_pmp_0_cfg_x; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_0_cfg_w = csr_io_pmp_0_cfg_w; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_0_cfg_r = csr_io_pmp_0_cfg_r; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_0_addr = csr_io_pmp_0_addr; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_0_mask = csr_io_pmp_0_mask; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_1_cfg_l = csr_io_pmp_1_cfg_l; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_1_cfg_a = csr_io_pmp_1_cfg_a; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_1_cfg_x = csr_io_pmp_1_cfg_x; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_1_cfg_w = csr_io_pmp_1_cfg_w; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_1_cfg_r = csr_io_pmp_1_cfg_r; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_1_addr = csr_io_pmp_1_addr; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_1_mask = csr_io_pmp_1_mask; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_2_cfg_l = csr_io_pmp_2_cfg_l; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_2_cfg_a = csr_io_pmp_2_cfg_a; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_2_cfg_x = csr_io_pmp_2_cfg_x; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_2_cfg_w = csr_io_pmp_2_cfg_w; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_2_cfg_r = csr_io_pmp_2_cfg_r; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_2_addr = csr_io_pmp_2_addr; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_2_mask = csr_io_pmp_2_mask; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_3_cfg_l = csr_io_pmp_3_cfg_l; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_3_cfg_a = csr_io_pmp_3_cfg_a; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_3_cfg_x = csr_io_pmp_3_cfg_x; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_3_cfg_w = csr_io_pmp_3_cfg_w; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_3_cfg_r = csr_io_pmp_3_cfg_r; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_3_addr = csr_io_pmp_3_addr; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_3_mask = csr_io_pmp_3_mask; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_4_cfg_l = csr_io_pmp_4_cfg_l; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_4_cfg_a = csr_io_pmp_4_cfg_a; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_4_cfg_x = csr_io_pmp_4_cfg_x; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_4_cfg_w = csr_io_pmp_4_cfg_w; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_4_cfg_r = csr_io_pmp_4_cfg_r; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_4_addr = csr_io_pmp_4_addr; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_4_mask = csr_io_pmp_4_mask; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_5_cfg_l = csr_io_pmp_5_cfg_l; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_5_cfg_a = csr_io_pmp_5_cfg_a; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_5_cfg_x = csr_io_pmp_5_cfg_x; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_5_cfg_w = csr_io_pmp_5_cfg_w; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_5_cfg_r = csr_io_pmp_5_cfg_r; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_5_addr = csr_io_pmp_5_addr; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_5_mask = csr_io_pmp_5_mask; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_6_cfg_l = csr_io_pmp_6_cfg_l; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_6_cfg_a = csr_io_pmp_6_cfg_a; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_6_cfg_x = csr_io_pmp_6_cfg_x; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_6_cfg_w = csr_io_pmp_6_cfg_w; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_6_cfg_r = csr_io_pmp_6_cfg_r; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_6_addr = csr_io_pmp_6_addr; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_6_mask = csr_io_pmp_6_mask; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_7_cfg_l = csr_io_pmp_7_cfg_l; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_7_cfg_a = csr_io_pmp_7_cfg_a; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_7_cfg_x = csr_io_pmp_7_cfg_x; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_7_cfg_w = csr_io_pmp_7_cfg_w; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_7_cfg_r = csr_io_pmp_7_cfg_r; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_7_addr = csr_io_pmp_7_addr; // @[RocketCore.scala 696:14]
  assign io_ptw_pmp_7_mask = csr_io_pmp_7_mask; // @[RocketCore.scala 696:14]
  assign io_ptw_customCSRs_csrs_0_value = csr_io_customCSRs_0_value; // @[RocketCore.scala 694:79]
  assign io_fpu_inst = ibuf_io_inst_0_bits_inst_bits; // @[RocketCore.scala 820:15]
  assign io_fpu_fromint_data = ex_reg_rs_bypass_0 ? _T_1015 : _T_1016; // @[RocketCore.scala 821:23]
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm; // @[RocketCore.scala 682:18]
  assign io_fpu_dmem_resp_val = dmem_resp_valid & io_dmem_resp_bits_tag[0]; // @[RocketCore.scala 822:24]
  assign io_fpu_dmem_resp_type = {{1'd0}, io_dmem_resp_bits_size}; // @[RocketCore.scala 824:25]
  assign io_fpu_dmem_resp_tag = io_dmem_resp_bits_tag[5:1]; // @[RocketCore.scala 825:24]
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data_word_bypass; // @[RocketCore.scala 823:25]
  assign io_fpu_valid = ~ctrl_killd & id_ctrl_fp; // @[RocketCore.scala 817:16]
  assign io_fpu_killx = _T_1157 | ~ex_reg_valid; // @[RocketCore.scala 818:16]
  assign io_fpu_killm = _T_1442 | ~mem_reg_valid; // @[RocketCore.scala 819:16]
  assign io_wfi = csr_io_status_wfi; // @[RocketCore.scala 855:10]
  assign ibuf_clock = clock;
  assign ibuf_reset = reset;
  assign ibuf_io_imem_valid = io_imem_resp_valid; // @[RocketCore.scala 252:16]
  assign ibuf_io_imem_bits_btb_taken = io_imem_resp_bits_btb_taken; // @[RocketCore.scala 252:16]
  assign ibuf_io_imem_bits_btb_bridx = io_imem_resp_bits_btb_bridx; // @[RocketCore.scala 252:16]
  assign ibuf_io_imem_bits_btb_entry = io_imem_resp_bits_btb_entry; // @[RocketCore.scala 252:16]
  assign ibuf_io_imem_bits_btb_bht_history = io_imem_resp_bits_btb_bht_history; // @[RocketCore.scala 252:16]
  assign ibuf_io_imem_bits_pc = io_imem_resp_bits_pc; // @[RocketCore.scala 252:16]
  assign ibuf_io_imem_bits_data = io_imem_resp_bits_data; // @[RocketCore.scala 252:16]
  assign ibuf_io_imem_bits_xcpt_pf_inst = io_imem_resp_bits_xcpt_pf_inst; // @[RocketCore.scala 252:16]
  assign ibuf_io_imem_bits_xcpt_ae_inst = io_imem_resp_bits_xcpt_ae_inst; // @[RocketCore.scala 252:16]
  assign ibuf_io_imem_bits_replay = io_imem_resp_bits_replay; // @[RocketCore.scala 252:16]
  assign ibuf_io_kill = take_pc_wb | take_pc_mem; // @[RocketCore.scala 253:16]
  assign ibuf_io_inst_0_ready = ~ctrl_stalld; // @[RocketCore.scala 796:25]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_ungated_clock = clock; // @[RocketCore.scala 674:24]
  assign csr_io_interrupts_debug = io_interrupts_debug; // @[RocketCore.scala 680:21]
  assign csr_io_interrupts_mtip = io_interrupts_mtip; // @[RocketCore.scala 680:21]
  assign csr_io_interrupts_msip = io_interrupts_msip; // @[RocketCore.scala 680:21]
  assign csr_io_interrupts_meip = io_interrupts_meip; // @[RocketCore.scala 680:21]
  assign csr_io_interrupts_seip = io_interrupts_seip; // @[RocketCore.scala 680:21]
  assign csr_io_hartid = io_hartid; // @[RocketCore.scala 681:17]
  assign csr_io_rw_addr = wb_reg_inst[31:20]; // @[RocketCore.scala 697:18]
  assign csr_io_rw_cmd = wb_ctrl_csr & ~_T_1565; // @[RocketCore.scala 698:17]
  assign csr_io_rw_wdata = wb_reg_wdata; // @[RocketCore.scala 699:19]
  assign csr_io_decode_0_csr = ibuf_io_inst_0_bits_raw[31:20]; // @[RocketCore.scala 675:24]
  assign csr_io_exception = _T_1481 | _T_1476; // @[RocketCore.scala 676:20]
  assign csr_io_retire = _T_1513 & ~wb_xcpt; // @[RocketCore.scala 678:17]
  assign csr_io_cause = wb_reg_xcpt ? wb_reg_cause : {{60'd0}, _T_1486}; // @[RocketCore.scala 677:16]
  assign csr_io_pc = wb_reg_pc; // @[RocketCore.scala 687:13]
  assign csr_io_tval = tval_valid ? _T_1562 : 40'h0; // @[RocketCore.scala 692:15]
  assign csr_io_fcsr_flags_valid = io_fpu_fcsr_flags_valid; // @[RocketCore.scala 683:21]
  assign csr_io_fcsr_flags_bits = io_fpu_fcsr_flags_bits; // @[RocketCore.scala 683:21]
  assign csr_io_inst_0 = {_T_1531,wb_reg_raw_inst[15:0]}; // @[RocketCore.scala 679:18]
  assign bpu_io_status_debug = csr_io_status_debug; // @[RocketCore.scala 318:17]
  assign bpu_io_status_prv = csr_io_status_prv; // @[RocketCore.scala 318:17]
  assign bpu_io_bp_0_control_action = csr_io_bp_0_control_action; // @[RocketCore.scala 319:13]
  assign bpu_io_bp_0_control_tmatch = csr_io_bp_0_control_tmatch; // @[RocketCore.scala 319:13]
  assign bpu_io_bp_0_control_m = csr_io_bp_0_control_m; // @[RocketCore.scala 319:13]
  assign bpu_io_bp_0_control_s = csr_io_bp_0_control_s; // @[RocketCore.scala 319:13]
  assign bpu_io_bp_0_control_u = csr_io_bp_0_control_u; // @[RocketCore.scala 319:13]
  assign bpu_io_bp_0_control_x = csr_io_bp_0_control_x; // @[RocketCore.scala 319:13]
  assign bpu_io_bp_0_control_w = csr_io_bp_0_control_w; // @[RocketCore.scala 319:13]
  assign bpu_io_bp_0_control_r = csr_io_bp_0_control_r; // @[RocketCore.scala 319:13]
  assign bpu_io_bp_0_address = csr_io_bp_0_address; // @[RocketCore.scala 319:13]
  assign bpu_io_pc = ibuf_io_pc[38:0]; // @[RocketCore.scala 320:13]
  assign bpu_io_ea = mem_reg_wdata[38:0]; // @[RocketCore.scala 321:13]
  assign alu_io_dw = ex_ctrl_alu_dw; // @[RocketCore.scala 378:13]
  assign alu_io_fn = ex_ctrl_alu_fn; // @[RocketCore.scala 379:13]
  assign alu_io_in2 = _T_1096 ? $signed({{60{_T_1091[3]}},_T_1091}) : $signed(_T_1095); // @[RocketCore.scala 380:14]
  assign alu_io_in1 = _T_1089 ? $signed({{24{ex_reg_pc[39]}},ex_reg_pc}) : $signed(_T_1088); // @[RocketCore.scala 381:14]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_req_valid = ex_reg_valid & ex_ctrl_div; // @[RocketCore.scala 402:20]
  assign div_io_req_bits_fn = ex_ctrl_alu_fn; // @[RocketCore.scala 404:22]
  assign div_io_req_bits_dw = ex_ctrl_alu_dw; // @[RocketCore.scala 403:22]
  assign div_io_req_bits_in1 = ex_reg_rs_bypass_0 ? _T_1015 : _T_1016; // @[RocketCore.scala 405:23]
  assign div_io_req_bits_in2 = ex_reg_rs_bypass_1 ? _T_1022 : _T_1023; // @[RocketCore.scala 406:23]
  assign div_io_req_bits_tag = ex_reg_inst[11:7]; // @[RocketCore.scala 407:23]
  assign div_io_kill = killm_common & _T_1445; // @[RocketCore.scala 580:15]
  assign div_io_resp_ready = _T_1511 ? 1'h0 : ~wb_wxd; // @[RocketCore.scala 641:21 RocketCore.scala 655:23]
  assign Rocket_cov_read_addr = Rocket_state;
  assign Rocket_cov_read_data = Rocket_cov[Rocket_cov_read_addr]; // @[Coverage map for Rocket]
  assign Rocket_cov_write_data = 1'h1;
  assign Rocket_cov_write_addr = Rocket_state;
  assign Rocket_cov_write_mask = 1'h1;
  assign Rocket_cov_write_en = 1'h1;
  assign mux_cond_0 = _T_1529;
  assign mux_cond_1 = _T_1557;
  assign mux_cond_2 = _T_1521;
  assign mux_cond_3 = _T_1309;
  assign mux_cond_4 = _T_1526;
  assign mux_cond_5 = _T_1525;
  assign mem_reg_slow_bypass_shl = {mem_reg_slow_bypass, 16'h0};
  assign mem_reg_slow_bypass_pad = {3'h0,mem_reg_slow_bypass_shl};
  assign ex_ctrl_sel_alu1_shl = ex_ctrl_sel_alu1;
  assign ex_ctrl_sel_alu1_pad = {18'h0,ex_ctrl_sel_alu1_shl};
  assign ex_ctrl_wxd_shl = {ex_ctrl_wxd, 2'h0};
  assign ex_ctrl_wxd_pad = {17'h0,ex_ctrl_wxd_shl};
  assign wb_ctrl_rxs2_shl = {wb_ctrl_rxs2, 18'h0};
  assign wb_ctrl_rxs2_pad = {1'h0,wb_ctrl_rxs2_shl};
  assign mem_reg_store_shl = {mem_reg_store, 16'h0};
  assign mem_reg_store_pad = {3'h0,mem_reg_store_shl};
  assign wb_reg_valid_shl = {wb_reg_valid, 6'h0};
  assign wb_reg_valid_pad = {13'h0,wb_reg_valid_shl};
  assign mem_ctrl_jal_shl = {mem_ctrl_jal, 2'h0};
  assign mem_ctrl_jal_pad = {17'h0,mem_ctrl_jal_shl};
  assign mem_br_taken_shl = {mem_br_taken, 16'h0};
  assign mem_br_taken_pad = {3'h0,mem_br_taken_shl};
  assign ex_ctrl_jalr_shl = {ex_ctrl_jalr, 13'h0};
  assign ex_ctrl_jalr_pad = {6'h0,ex_ctrl_jalr_shl};
  assign wb_ctrl_rfs2_shl = {wb_ctrl_rfs2, 11'h0};
  assign wb_ctrl_rfs2_pad = {8'h0,wb_ctrl_rfs2_shl};
  assign ex_ctrl_sel_imm_shl = {ex_ctrl_sel_imm, 7'h0};
  assign ex_ctrl_sel_imm_pad = {10'h0,ex_ctrl_sel_imm_shl};
  assign mem_ctrl_mem_shl = mem_ctrl_mem;
  assign mem_ctrl_mem_pad = {19'h0,mem_ctrl_mem_shl};
  assign wb_reg_xcpt_shl = {wb_reg_xcpt, 6'h0};
  assign wb_reg_xcpt_pad = {13'h0,wb_reg_xcpt_shl};
  assign ex_reg_xcpt_interrupt_shl = {ex_reg_xcpt_interrupt, 11'h0};
  assign ex_reg_xcpt_interrupt_pad = {8'h0,ex_reg_xcpt_interrupt_shl};
  assign mem_ctrl_branch_shl = {mem_ctrl_branch, 9'h0};
  assign mem_ctrl_branch_pad = {10'h0,mem_ctrl_branch_shl};
  assign ex_ctrl_fp_shl = ex_ctrl_fp;
  assign ex_ctrl_fp_pad = {19'h0,ex_ctrl_fp_shl};
  assign ex_reg_mem_size_shl = {ex_reg_mem_size, 8'h0};
  assign ex_reg_mem_size_pad = {10'h0,ex_reg_mem_size_shl};
  assign mem_ctrl_wfd_shl = {mem_ctrl_wfd, 1'h0};
  assign mem_ctrl_wfd_pad = {18'h0,mem_ctrl_wfd_shl};
  assign mem_reg_load_shl = {mem_reg_load, 18'h0};
  assign mem_reg_load_pad = {1'h0,mem_reg_load_shl};
  assign mem_reg_flush_pipe_shl = {mem_reg_flush_pipe, 18'h0};
  assign mem_reg_flush_pipe_pad = {1'h0,mem_reg_flush_pipe_shl};
  assign wb_reg_replay_shl = {wb_reg_replay, 11'h0};
  assign wb_reg_replay_pad = {8'h0,wb_reg_replay_shl};
  assign id_reg_pause_shl = {id_reg_pause, 8'h0};
  assign id_reg_pause_pad = {11'h0,id_reg_pause_shl};
  assign wb_ctrl_rxs1_shl = {wb_ctrl_rxs1, 3'h0};
  assign wb_ctrl_rxs1_pad = {16'h0,wb_ctrl_rxs1_shl};
  assign ex_ctrl_rxs2_shl = {ex_ctrl_rxs2, 17'h0};
  assign ex_ctrl_rxs2_pad = {2'h0,ex_ctrl_rxs2_shl};
  assign ex_reg_replay_shl = {ex_reg_replay, 1'h0};
  assign ex_reg_replay_pad = {18'h0,ex_reg_replay_shl};
  assign mem_ctrl_div_shl = {mem_ctrl_div, 7'h0};
  assign mem_ctrl_div_pad = {12'h0,mem_ctrl_div_shl};
  assign wb_ctrl_wfd_shl = {wb_ctrl_wfd, 12'h0};
  assign wb_ctrl_wfd_pad = {7'h0,wb_ctrl_wfd_shl};
  assign wb_ctrl_mem_shl = {wb_ctrl_mem, 12'h0};
  assign wb_ctrl_mem_pad = {7'h0,wb_ctrl_mem_shl};
  assign wb_reg_flush_pipe_shl = {wb_reg_flush_pipe, 19'h0};
  assign wb_reg_flush_pipe_pad = wb_reg_flush_pipe_shl;
  assign mem_reg_rvc_shl = {mem_reg_rvc, 8'h0};
  assign mem_reg_rvc_pad = {11'h0,mem_reg_rvc_shl};
  assign mem_reg_xcpt_interrupt_shl = {mem_reg_xcpt_interrupt, 8'h0};
  assign mem_reg_xcpt_interrupt_pad = {11'h0,mem_reg_xcpt_interrupt_shl};
  assign ex_ctrl_mem_shl = {ex_ctrl_mem, 3'h0};
  assign ex_ctrl_mem_pad = {16'h0,ex_ctrl_mem_shl};
  assign ex_ctrl_sel_alu2_shl = {ex_ctrl_sel_alu2, 9'h0};
  assign ex_ctrl_sel_alu2_pad = {9'h0,ex_ctrl_sel_alu2_shl};
  assign id_reg_fence_shl = {id_reg_fence, 4'h0};
  assign id_reg_fence_pad = {15'h0,id_reg_fence_shl};
  assign mem_ctrl_wxd_shl = {mem_ctrl_wxd, 14'h0};
  assign mem_ctrl_wxd_pad = {5'h0,mem_ctrl_wxd_shl};
  assign mem_reg_xcpt_shl = {mem_reg_xcpt, 2'h0};
  assign mem_reg_xcpt_pad = {17'h0,mem_reg_xcpt_shl};
  assign ex_reg_valid_shl = {ex_reg_valid, 19'h0};
  assign ex_reg_valid_pad = ex_reg_valid_shl;
  assign ex_ctrl_div_shl = {ex_ctrl_div, 14'h0};
  assign ex_ctrl_div_pad = {5'h0,ex_ctrl_div_shl};
  assign ex_ctrl_wfd_shl = {ex_ctrl_wfd, 5'h0};
  assign ex_ctrl_wfd_pad = {14'h0,ex_ctrl_wfd_shl};
  assign wb_ctrl_rfs1_shl = {wb_ctrl_rfs1, 4'h0};
  assign wb_ctrl_rfs1_pad = {15'h0,wb_ctrl_rfs1_shl};
  assign mem_ctrl_fp_shl = {mem_ctrl_fp, 7'h0};
  assign mem_ctrl_fp_pad = {12'h0,mem_ctrl_fp_shl};
  assign mem_reg_sfence_shl = {mem_reg_sfence, 11'h0};
  assign mem_reg_sfence_pad = {8'h0,mem_reg_sfence_shl};
  assign wb_ctrl_div_shl = {wb_ctrl_div, 12'h0};
  assign wb_ctrl_div_pad = {7'h0,wb_ctrl_div_shl};
  assign mem_reg_replay_shl = {mem_reg_replay, 9'h0};
  assign mem_reg_replay_pad = {10'h0,mem_reg_replay_shl};
  assign ex_reg_rvc_shl = {ex_reg_rvc, 14'h0};
  assign ex_reg_rvc_pad = {5'h0,ex_reg_rvc_shl};
  assign blocked_shl = {blocked, 6'h0};
  assign blocked_pad = {13'h0,blocked_shl};
  assign mem_reg_valid_shl = {mem_reg_valid, 5'h0};
  assign mem_reg_valid_pad = {14'h0,mem_reg_valid_shl};
  assign mem_ctrl_jalr_shl = {mem_ctrl_jalr, 16'h0};
  assign mem_ctrl_jalr_pad = {3'h0,mem_ctrl_jalr_shl};
  assign wb_ctrl_wxd_shl = {wb_ctrl_wxd, 8'h0};
  assign wb_ctrl_wxd_pad = {11'h0,wb_ctrl_wxd_shl};
  assign mux_cond_0_shl = {mux_cond_0, 17'h0};
  assign mux_cond_0_pad = {2'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 17'h0};
  assign mux_cond_1_pad = {2'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 9'h0};
  assign mux_cond_2_pad = {10'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 10'h0};
  assign mux_cond_3_pad = {9'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 15'h0};
  assign mux_cond_4_pad = {4'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = mux_cond_5;
  assign mux_cond_5_pad = {19'h0,mux_cond_5_shl};
  assign ex_reg_rs_lsb_0_shl = {ex_reg_rs_lsb_0, 9'h0};
  assign ex_reg_rs_lsb_0_pad = {9'h0,ex_reg_rs_lsb_0_shl};
  assign ex_reg_rs_lsb_1_shl = {ex_reg_rs_lsb_1, 9'h0};
  assign ex_reg_rs_lsb_1_pad = {9'h0,ex_reg_rs_lsb_1_shl};
  assign ex_reg_rs_bypass_0_shl = {ex_reg_rs_bypass_0, 13'h0};
  assign ex_reg_rs_bypass_0_pad = {6'h0,ex_reg_rs_bypass_0_shl};
  assign ex_reg_rs_bypass_1_shl = {ex_reg_rs_bypass_1, 13'h0};
  assign ex_reg_rs_bypass_1_pad = {6'h0,ex_reg_rs_bypass_1_shl};
  assign Rocket_xor32 = ex_ctrl_sel_alu1_pad ^ ex_ctrl_wxd_pad;
  assign Rocket_xor15 = mem_reg_slow_bypass_pad ^ Rocket_xor32;
  assign Rocket_xor33 = wb_ctrl_rxs2_pad ^ mem_reg_store_pad;
  assign Rocket_xor34 = wb_reg_valid_pad ^ mem_ctrl_jal_pad;
  assign Rocket_xor16 = Rocket_xor33 ^ Rocket_xor34;
  assign Rocket_xor7 = Rocket_xor15 ^ Rocket_xor16;
  assign Rocket_xor36 = ex_ctrl_jalr_pad ^ wb_ctrl_rfs2_pad;
  assign Rocket_xor17 = mem_br_taken_pad ^ Rocket_xor36;
  assign Rocket_xor37 = ex_ctrl_sel_imm_pad ^ mem_ctrl_mem_pad;
  assign Rocket_xor38 = wb_reg_xcpt_pad ^ ex_reg_xcpt_interrupt_pad;
  assign Rocket_xor18 = Rocket_xor37 ^ Rocket_xor38;
  assign Rocket_xor8 = Rocket_xor17 ^ Rocket_xor18;
  assign Rocket_xor3 = Rocket_xor7 ^ Rocket_xor8;
  assign Rocket_xor40 = ex_ctrl_fp_pad ^ ex_reg_mem_size_pad;
  assign Rocket_xor19 = mem_ctrl_branch_pad ^ Rocket_xor40;
  assign Rocket_xor41 = mem_ctrl_wfd_pad ^ mem_reg_load_pad;
  assign Rocket_xor42 = mem_reg_flush_pipe_pad ^ wb_reg_replay_pad;
  assign Rocket_xor20 = Rocket_xor41 ^ Rocket_xor42;
  assign Rocket_xor9 = Rocket_xor19 ^ Rocket_xor20;
  assign Rocket_xor43 = id_reg_pause_pad ^ wb_ctrl_rxs1_pad;
  assign Rocket_xor44 = ex_ctrl_rxs2_pad ^ ex_reg_replay_pad;
  assign Rocket_xor21 = Rocket_xor43 ^ Rocket_xor44;
  assign Rocket_xor45 = mem_ctrl_div_pad ^ wb_ctrl_wfd_pad;
  assign Rocket_xor46 = wb_ctrl_mem_pad ^ wb_reg_flush_pipe_pad;
  assign Rocket_xor22 = Rocket_xor45 ^ Rocket_xor46;
  assign Rocket_xor10 = Rocket_xor21 ^ Rocket_xor22;
  assign Rocket_xor4 = Rocket_xor9 ^ Rocket_xor10;
  assign Rocket_xor1 = Rocket_xor3 ^ Rocket_xor4;
  assign Rocket_xor48 = mem_reg_xcpt_interrupt_pad ^ ex_ctrl_mem_pad;
  assign Rocket_xor23 = mem_reg_rvc_pad ^ Rocket_xor48;
  assign Rocket_xor49 = ex_ctrl_sel_alu2_pad ^ id_reg_fence_pad;
  assign Rocket_xor50 = mem_ctrl_wxd_pad ^ mem_reg_xcpt_pad;
  assign Rocket_xor24 = Rocket_xor49 ^ Rocket_xor50;
  assign Rocket_xor11 = Rocket_xor23 ^ Rocket_xor24;
  assign Rocket_xor51 = ex_reg_valid_pad ^ ex_ctrl_div_pad;
  assign Rocket_xor52 = ex_ctrl_wfd_pad ^ wb_ctrl_rfs1_pad;
  assign Rocket_xor25 = Rocket_xor51 ^ Rocket_xor52;
  assign Rocket_xor53 = mem_ctrl_fp_pad ^ mem_reg_sfence_pad;
  assign Rocket_xor54 = wb_ctrl_div_pad ^ mem_reg_replay_pad;
  assign Rocket_xor26 = Rocket_xor53 ^ Rocket_xor54;
  assign Rocket_xor12 = Rocket_xor25 ^ Rocket_xor26;
  assign Rocket_xor5 = Rocket_xor11 ^ Rocket_xor12;
  assign Rocket_xor56 = blocked_pad ^ mem_reg_valid_pad;
  assign Rocket_xor27 = ex_reg_rvc_pad ^ Rocket_xor56;
  assign Rocket_xor57 = mem_ctrl_jalr_pad ^ wb_ctrl_wxd_pad;
  assign Rocket_xor58 = mux_cond_0_pad ^ mux_cond_1_pad;
  assign Rocket_xor28 = Rocket_xor57 ^ Rocket_xor58;
  assign Rocket_xor13 = Rocket_xor27 ^ Rocket_xor28;
  assign Rocket_xor59 = mux_cond_2_pad ^ mux_cond_3_pad;
  assign Rocket_xor60 = mux_cond_4_pad ^ mux_cond_5_pad;
  assign Rocket_xor29 = Rocket_xor59 ^ Rocket_xor60;
  assign Rocket_xor61 = ex_reg_rs_lsb_0_pad ^ ex_reg_rs_lsb_1_pad;
  assign Rocket_xor62 = ex_reg_rs_bypass_0_pad ^ ex_reg_rs_bypass_1_pad;
  assign Rocket_xor30 = Rocket_xor61 ^ Rocket_xor62;
  assign Rocket_xor14 = Rocket_xor29 ^ Rocket_xor30;
  assign Rocket_xor6 = Rocket_xor13 ^ Rocket_xor14;
  assign Rocket_xor2 = Rocket_xor5 ^ Rocket_xor6;
  assign Rocket_xor0 = Rocket_xor1 ^ Rocket_xor2;
  assign alu_sum = Rocket_covSum + alu_io_covSum;
  assign csr_sum = alu_sum + csr_io_covSum;
  assign div_sum = csr_sum + div_io_covSum;
  assign bpu_sum = div_sum + bpu_io_covSum;
  assign ibuf_sum = bpu_sum + ibuf_io_covSum;
  assign PlusArgTimeout_sum = ibuf_sum + PlusArgTimeout_io_covSum;
  assign io_covSum = PlusArgTimeout_sum;
  assign alu_metaAssert_wire = alu_metaAssert;
  assign bpu_metaAssert_wire = bpu_metaAssert;
  assign csr_metaAssert_wire = csr_metaAssert;
  assign ibuf_metaAssert_wire = ibuf_metaAssert;
  assign PlusArgTimeout_metaAssert_wire = PlusArgTimeout_metaAssert;
  assign div_metaAssert_wire = div_metaAssert;
  assign Rocket_or4 = alu_metaAssert_wire | PlusArgTimeout_metaAssert_wire;
  assign Rocket_or1 = ibuf_metaAssert_wire | Rocket_or4;
  assign Rocket_or6 = div_metaAssert_wire | csr_metaAssert_wire;
  assign Rocket_or2 = bpu_metaAssert_wire | Rocket_or6;
  assign Rocket_or0 = Rocket_or1 | Rocket_or2;
  assign metaAssert = Rocket_metaAssert;
  assign csr_metaReset = metaReset | csr_halt;
  assign div_metaReset = metaReset | div_halt;
  assign ibuf_metaReset = metaReset | ibuf_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 31; initvar = initvar+1)
    _T_815[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  _RAND_2 = {2{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  id_reg_pause = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  imem_might_request_reg = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ex_ctrl_fp = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ex_ctrl_branch = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ex_ctrl_jal = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ex_ctrl_jalr = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  ex_ctrl_rxs2 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  ex_ctrl_rxs1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  ex_ctrl_sel_alu2 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  ex_ctrl_sel_alu1 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  ex_ctrl_sel_imm = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  ex_ctrl_alu_dw = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  ex_ctrl_alu_fn = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  ex_ctrl_mem = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  ex_ctrl_mem_cmd = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  ex_ctrl_rfs1 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  ex_ctrl_rfs2 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  ex_ctrl_wfd = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  ex_ctrl_div = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  ex_ctrl_wxd = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  ex_ctrl_csr = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  ex_ctrl_fence_i = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  mem_ctrl_fp = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mem_ctrl_branch = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mem_ctrl_jal = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  mem_ctrl_jalr = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  mem_ctrl_rxs2 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  mem_ctrl_rxs1 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  mem_ctrl_mem = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  mem_ctrl_rfs1 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  mem_ctrl_rfs2 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  mem_ctrl_wfd = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  mem_ctrl_div = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  mem_ctrl_wxd = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  mem_ctrl_csr = _RAND_37[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  mem_ctrl_fence_i = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  wb_ctrl_rxs2 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  wb_ctrl_rxs1 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  wb_ctrl_mem = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  wb_ctrl_rfs1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  wb_ctrl_rfs2 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  wb_ctrl_wfd = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  wb_ctrl_div = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  wb_ctrl_wxd = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  wb_ctrl_csr = _RAND_47[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  wb_ctrl_fence_i = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  ex_reg_xcpt_interrupt = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  ex_reg_valid = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  ex_reg_rvc = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  ex_reg_btb_resp_entry = _RAND_52[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  ex_reg_btb_resp_bht_history = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  ex_reg_xcpt = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  ex_reg_flush_pipe = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  ex_reg_load_use = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  ex_reg_cause = _RAND_57[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  ex_reg_replay = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {2{`RANDOM}};
  ex_reg_pc = _RAND_59[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  ex_reg_mem_size = _RAND_60[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  ex_reg_inst = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  ex_reg_raw_inst = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  mem_reg_xcpt_interrupt = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  mem_reg_valid = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  mem_reg_rvc = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  mem_reg_btb_resp_entry = _RAND_66[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  mem_reg_btb_resp_bht_history = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  mem_reg_xcpt = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  mem_reg_replay = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  mem_reg_flush_pipe = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {2{`RANDOM}};
  mem_reg_cause = _RAND_71[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  mem_reg_slow_bypass = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  mem_reg_load = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  mem_reg_store = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  mem_reg_sfence = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{`RANDOM}};
  mem_reg_pc = _RAND_76[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  mem_reg_inst = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  mem_reg_mem_size = _RAND_78[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  mem_reg_raw_inst = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {2{`RANDOM}};
  mem_reg_wdata = _RAND_80[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {2{`RANDOM}};
  mem_reg_rs2 = _RAND_81[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  mem_br_taken = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  wb_reg_valid = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  wb_reg_xcpt = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  wb_reg_replay = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  wb_reg_flush_pipe = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {2{`RANDOM}};
  wb_reg_cause = _RAND_87[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  wb_reg_sfence = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {2{`RANDOM}};
  wb_reg_pc = _RAND_89[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  wb_reg_mem_size = _RAND_90[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  wb_reg_inst = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  wb_reg_raw_inst = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {2{`RANDOM}};
  wb_reg_wdata = _RAND_93[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  id_reg_fence = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  ex_reg_rs_bypass_0 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  ex_reg_rs_bypass_1 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  ex_reg_rs_lsb_0 = _RAND_97[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  ex_reg_rs_lsb_1 = _RAND_98[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {2{`RANDOM}};
  ex_reg_rs_msb_0 = _RAND_99[61:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {2{`RANDOM}};
  ex_reg_rs_msb_1 = _RAND_100[61:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_1574 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_1687 = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  blocked = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_1445 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {2{`RANDOM}};
  _T_1866 = _RAND_105[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {2{`RANDOM}};
  coreMonitorBundle_rd0val = _RAND_106[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {2{`RANDOM}};
  _T_1869 = _RAND_107[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {2{`RANDOM}};
  coreMonitorBundle_rd1val = _RAND_108[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  Rocket_state = _RAND_109[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    Rocket_cov[initvar] = _RAND_110[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  Rocket_covSum = _RAND_111[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  Rocket_metaAssert = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_815__T_1524_en & _T_815__T_1524_mask) begin
      _T_815[_T_815__T_1524_addr] <= _T_815__T_1524_data; // @[RocketCore.scala 1014:15]
    end
    if (metaReset) begin
      id_reg_pause <= 1'h0;
    end else if (unpause) begin
      id_reg_pause <= 1'h0;
    end else if (~ctrl_killd) begin
      id_reg_pause <= _GEN_1;
    end
    if (metaReset) begin
      imem_might_request_reg <= 1'h0;
    end else begin
      imem_might_request_reg <= _T_1774 | io_ptw_customCSRs_csrs_0_value[1];
    end
    if (metaReset) begin
      ex_ctrl_fp <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_fp <= id_ctrl_fp;
    end
    if (metaReset) begin
      ex_ctrl_branch <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_branch <= id_ctrl_branch;
    end
    if (metaReset) begin
      ex_ctrl_jal <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_jal <= id_ctrl_jal;
    end
    if (metaReset) begin
      ex_ctrl_jalr <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_jalr <= id_ctrl_jalr;
    end
    if (metaReset) begin
      ex_ctrl_rxs2 <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_rxs2 <= id_ctrl_rxs2;
    end
    if (metaReset) begin
      ex_ctrl_rxs1 <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_rxs1 <= id_ctrl_rxs1;
    end
    if (metaReset) begin
      ex_ctrl_sel_alu2 <= 2'h0;
    end else if (~ctrl_killd) begin
      if (id_xcpt) begin
        if (_T_1118) begin
          ex_ctrl_sel_alu2 <= 2'h0;
        end else if (_T_1115) begin
          ex_ctrl_sel_alu2 <= 2'h1;
        end else begin
          ex_ctrl_sel_alu2 <= 2'h0;
        end
      end else begin
        ex_ctrl_sel_alu2 <= id_ctrl_sel_alu2;
      end
    end
    if (metaReset) begin
      ex_ctrl_sel_alu1 <= 2'h0;
    end else if (~ctrl_killd) begin
      if (id_xcpt) begin
        if (_T_1118) begin
          ex_ctrl_sel_alu1 <= 2'h2;
        end else if (_T_1115) begin
          ex_ctrl_sel_alu1 <= 2'h2;
        end else begin
          ex_ctrl_sel_alu1 <= 2'h1;
        end
      end else begin
        ex_ctrl_sel_alu1 <= id_ctrl_sel_alu1;
      end
    end
    if (metaReset) begin
      ex_ctrl_sel_imm <= 3'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_sel_imm <= id_ctrl_sel_imm;
    end
    if (metaReset) begin
      ex_ctrl_alu_dw <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_alu_dw <= _GEN_9;
    end
    if (metaReset) begin
      ex_ctrl_alu_fn <= 4'h0;
    end else if (~ctrl_killd) begin
      if (id_xcpt) begin
        ex_ctrl_alu_fn <= 4'h0;
      end else begin
        ex_ctrl_alu_fn <= id_ctrl_alu_fn;
      end
    end
    if (metaReset) begin
      ex_ctrl_mem <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_mem <= id_ctrl_mem;
    end
    if (metaReset) begin
      ex_ctrl_mem_cmd <= 5'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_mem_cmd <= id_ctrl_mem_cmd;
    end
    if (metaReset) begin
      ex_ctrl_rfs1 <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_rfs1 <= id_ctrl_rfs1;
    end
    if (metaReset) begin
      ex_ctrl_rfs2 <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_rfs2 <= id_ctrl_rfs2;
    end
    if (metaReset) begin
      ex_ctrl_wfd <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_wfd <= id_ctrl_wfd;
    end
    if (metaReset) begin
      ex_ctrl_div <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_div <= id_ctrl_div;
    end
    if (metaReset) begin
      ex_ctrl_wxd <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_wxd <= id_ctrl_wxd;
    end
    if (metaReset) begin
      ex_ctrl_csr <= 3'h0;
    end else if (~ctrl_killd) begin
      if (id_csr_ren) begin
        ex_ctrl_csr <= 3'h2;
      end else begin
        ex_ctrl_csr <= id_ctrl_csr;
      end
    end
    if (metaReset) begin
      ex_ctrl_fence_i <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_fence_i <= id_ctrl_fence_i;
    end
    if (metaReset) begin
      mem_ctrl_fp <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_fp <= ex_ctrl_fp;
      end
    end
    if (metaReset) begin
      mem_ctrl_branch <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_branch <= ex_ctrl_branch;
      end
    end
    if (metaReset) begin
      mem_ctrl_jal <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_jal <= ex_ctrl_jal;
      end
    end
    if (metaReset) begin
      mem_ctrl_jalr <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_jalr <= ex_ctrl_jalr;
      end
    end
    if (metaReset) begin
      mem_ctrl_rxs2 <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_rxs2 <= ex_ctrl_rxs2;
      end
    end
    if (metaReset) begin
      mem_ctrl_rxs1 <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_rxs1 <= ex_ctrl_rxs1;
      end
    end
    if (metaReset) begin
      mem_ctrl_mem <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_mem <= ex_ctrl_mem;
      end
    end
    if (metaReset) begin
      mem_ctrl_rfs1 <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_rfs1 <= ex_ctrl_rfs1;
      end
    end
    if (metaReset) begin
      mem_ctrl_rfs2 <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_rfs2 <= ex_ctrl_rfs2;
      end
    end
    if (metaReset) begin
      mem_ctrl_wfd <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_wfd <= ex_ctrl_wfd;
      end
    end
    if (metaReset) begin
      mem_ctrl_div <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_div <= ex_ctrl_div;
      end
    end
    if (metaReset) begin
      mem_ctrl_wxd <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_wxd <= ex_ctrl_wxd;
      end
    end
    if (metaReset) begin
      mem_ctrl_csr <= 3'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_csr <= ex_ctrl_csr;
      end
    end
    if (metaReset) begin
      mem_ctrl_fence_i <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_ctrl_fence_i <= _GEN_77;
      end
    end
    if (metaReset) begin
      wb_ctrl_rxs2 <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_rxs2 <= mem_ctrl_rxs2;
    end
    if (metaReset) begin
      wb_ctrl_rxs1 <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_rxs1 <= mem_ctrl_rxs1;
    end
    if (metaReset) begin
      wb_ctrl_mem <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_mem <= mem_ctrl_mem;
    end
    if (metaReset) begin
      wb_ctrl_rfs1 <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_rfs1 <= mem_ctrl_rfs1;
    end
    if (metaReset) begin
      wb_ctrl_rfs2 <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_rfs2 <= mem_ctrl_rfs2;
    end
    if (metaReset) begin
      wb_ctrl_wfd <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_wfd <= mem_ctrl_wfd;
    end
    if (metaReset) begin
      wb_ctrl_div <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_div <= mem_ctrl_div;
    end
    if (metaReset) begin
      wb_ctrl_wxd <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_wxd <= mem_ctrl_wxd;
    end
    if (metaReset) begin
      wb_ctrl_csr <= 3'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_csr <= mem_ctrl_csr;
    end
    if (metaReset) begin
      wb_ctrl_fence_i <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_fence_i <= mem_ctrl_fence_i;
    end
    if (metaReset) begin
      ex_reg_xcpt_interrupt <= 1'h0;
    end else begin
      ex_reg_xcpt_interrupt <= _T_1102 & csr_io_interrupt;
    end
    if (metaReset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= ~ctrl_killd;
    end
    if (metaReset) begin
      ex_reg_rvc <= 1'h0;
    end else if (~ctrl_killd) begin
      if (id_xcpt) begin
        ex_reg_rvc <= _GEN_5;
      end else begin
        ex_reg_rvc <= ibuf_io_inst_0_bits_rvc;
      end
    end
    if (metaReset) begin
      ex_reg_btb_resp_entry <= 5'h0;
    end else if (_T_1148) begin
      ex_reg_btb_resp_entry <= ibuf_io_btb_resp_entry;
    end
    if (metaReset) begin
      ex_reg_btb_resp_bht_history <= 8'h0;
    end else if (_T_1148) begin
      ex_reg_btb_resp_bht_history <= ibuf_io_btb_resp_bht_history;
    end
    if (metaReset) begin
      ex_reg_xcpt <= 1'h0;
    end else begin
      ex_reg_xcpt <= ~ctrl_killd & id_xcpt;
    end
    if (metaReset) begin
      ex_reg_flush_pipe <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_reg_flush_pipe <= _T_1119;
    end
    if (metaReset) begin
      ex_reg_load_use <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_reg_load_use <= id_load_use;
    end
    if (metaReset) begin
      ex_reg_cause <= 64'h0;
    end else if (_T_1148) begin
      if (csr_io_interrupt) begin
        ex_reg_cause <= csr_io_interrupt_cause;
      end else begin
        ex_reg_cause <= {{60'd0}, _T_983};
      end
    end
    if (metaReset) begin
      ex_reg_replay <= 1'h0;
    end else begin
      ex_reg_replay <= _T_1102 & ibuf_io_inst_0_bits_replay;
    end
    if (metaReset) begin
      ex_reg_pc <= 40'h0;
    end else if (_T_1148) begin
      ex_reg_pc <= ibuf_io_pc;
    end
    if (metaReset) begin
      ex_reg_mem_size <= 2'h0;
    end else if (~ctrl_killd) begin
      if (_T_1123) begin
        ex_reg_mem_size <= _T_1126;
      end else begin
        ex_reg_mem_size <= ibuf_io_inst_0_bits_inst_bits[13:12];
      end
    end
    if (metaReset) begin
      ex_reg_inst <= 32'h0;
    end else if (_T_1148) begin
      ex_reg_inst <= ibuf_io_inst_0_bits_inst_bits;
    end
    if (metaReset) begin
      ex_reg_raw_inst <= 32'h0;
    end else if (_T_1148) begin
      ex_reg_raw_inst <= ibuf_io_inst_0_bits_raw;
    end
    if (metaReset) begin
      mem_reg_xcpt_interrupt <= 1'h0;
    end else begin
      mem_reg_xcpt_interrupt <= ~take_pc_mem_wb & ex_reg_xcpt_interrupt;
    end
    if (metaReset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= ~ctrl_killx;
    end
    if (metaReset) begin
      mem_reg_rvc <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_rvc <= ex_reg_rvc;
      end
    end
    if (metaReset) begin
      mem_reg_btb_resp_entry <= 5'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
      end
    end
    if (metaReset) begin
      mem_reg_btb_resp_bht_history <= 8'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
      end
    end
    if (metaReset) begin
      mem_reg_xcpt <= 1'h0;
    end else begin
      mem_reg_xcpt <= ~ctrl_killx & ex_xcpt;
    end
    if (metaReset) begin
      mem_reg_replay <= 1'h0;
    end else begin
      mem_reg_replay <= ~take_pc_mem_wb & replay_ex;
    end
    if (metaReset) begin
      mem_reg_flush_pipe <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_flush_pipe <= _GEN_78;
      end
    end
    if (metaReset) begin
      mem_reg_cause <= 64'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_cause <= ex_reg_cause;
      end
    end
    if (metaReset) begin
      mem_reg_slow_bypass <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_slow_bypass <= ex_slow_bypass;
      end
    end
    if (metaReset) begin
      mem_reg_load <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_load <= _T_1371;
      end
    end
    if (metaReset) begin
      mem_reg_store <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_store <= _T_1395;
      end
    end
    if (metaReset) begin
      mem_reg_sfence <= 1'h0;
    end else if (_T_1347) begin
      mem_reg_sfence <= 1'h0;
    end else if (ex_pc_valid) begin
      mem_reg_sfence <= ex_sfence;
    end
    if (metaReset) begin
      mem_reg_pc <= 40'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_pc <= ex_reg_pc;
      end
    end
    if (metaReset) begin
      mem_reg_inst <= 32'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_inst <= ex_reg_inst;
      end
    end
    if (metaReset) begin
      mem_reg_mem_size <= 2'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_mem_size <= ex_reg_mem_size;
      end
    end
    if (metaReset) begin
      mem_reg_raw_inst <= 32'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_raw_inst <= ex_reg_raw_inst;
      end
    end
    if (metaReset) begin
      mem_reg_wdata <= 64'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_reg_wdata <= _T_1396;
      end
    end
    if (metaReset) begin
      mem_reg_rs2 <= 64'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        if (_T_1399) begin
          if (_T_1401) begin
            mem_reg_rs2 <= _T_1405;
          end else if (_T_1406) begin
            mem_reg_rs2 <= _T_1409;
          end else if (_T_1410) begin
            mem_reg_rs2 <= _T_1412;
          end else if (ex_reg_rs_bypass_1) begin
            if (_T_1021) begin
              mem_reg_rs2 <= io_dmem_resp_bits_data_word_bypass;
            end else if (_T_1019) begin
              mem_reg_rs2 <= wb_reg_wdata;
            end else if (_T_1017) begin
              mem_reg_rs2 <= mem_reg_wdata;
            end else begin
              mem_reg_rs2 <= 64'h0;
            end
          end else begin
            mem_reg_rs2 <= _T_1023;
          end
        end
      end
    end
    if (metaReset) begin
      mem_br_taken <= 1'h0;
    end else if (!(_T_1347)) begin
      if (ex_pc_valid) begin
        mem_br_taken <= alu_io_cmp_out;
      end
    end
    if (metaReset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= ~ctrl_killm;
    end
    if (metaReset) begin
      wb_reg_xcpt <= 1'h0;
    end else begin
      wb_reg_xcpt <= mem_xcpt & ~take_pc_wb;
    end
    if (metaReset) begin
      wb_reg_replay <= 1'h0;
    end else begin
      wb_reg_replay <= replay_mem & ~take_pc_wb;
    end
    if (metaReset) begin
      wb_reg_flush_pipe <= 1'h0;
    end else begin
      wb_reg_flush_pipe <= ~ctrl_killm & mem_reg_flush_pipe;
    end
    if (metaReset) begin
      wb_reg_cause <= 64'h0;
    end else if (mem_pc_valid) begin
      if (_T_1421) begin
        wb_reg_cause <= mem_reg_cause;
      end else begin
        wb_reg_cause <= {{60'd0}, _T_1425};
      end
    end
    if (metaReset) begin
      wb_reg_sfence <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_reg_sfence <= mem_reg_sfence;
    end
    if (metaReset) begin
      wb_reg_pc <= 40'h0;
    end else if (mem_pc_valid) begin
      wb_reg_pc <= mem_reg_pc;
    end
    if (metaReset) begin
      wb_reg_mem_size <= 2'h0;
    end else if (mem_pc_valid) begin
      wb_reg_mem_size <= mem_reg_mem_size;
    end
    if (metaReset) begin
      wb_reg_inst <= 32'h0;
    end else if (mem_pc_valid) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if (metaReset) begin
      wb_reg_raw_inst <= 32'h0;
    end else if (mem_pc_valid) begin
      wb_reg_raw_inst <= mem_reg_raw_inst;
    end
    if (metaReset) begin
      wb_reg_wdata <= 64'h0;
    end else if (mem_pc_valid) begin
      if (_T_1457) begin
        wb_reg_wdata <= io_fpu_toint_data;
      end else begin
        wb_reg_wdata <= mem_int_wdata;
      end
    end
    if (metaReset) begin
      id_reg_fence <= 1'h0;
    end else if (reset) begin
      id_reg_fence <= 1'h0;
    end else if (~ctrl_killd) begin
      id_reg_fence <= _GEN_2;
    end else if (~id_mem_busy) begin
      id_reg_fence <= 1'h0;
    end
    if (metaReset) begin
      ex_reg_rs_bypass_0 <= 1'h0;
    end else if (~ctrl_killd) begin
      if (id_illegal_insn) begin
        ex_reg_rs_bypass_0 <= 1'h0;
      end else begin
        ex_reg_rs_bypass_0 <= do_bypass;
      end
    end
    if (metaReset) begin
      ex_reg_rs_bypass_1 <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_reg_rs_bypass_1 <= do_bypass_1;
    end
    if (metaReset) begin
      ex_reg_rs_lsb_0 <= 2'h0;
    end else if (~ctrl_killd) begin
      if (id_illegal_insn) begin
        ex_reg_rs_lsb_0 <= inst[1:0];
      end else if (_T_1132) begin
        ex_reg_rs_lsb_0 <= id_rs_0[1:0];
      end else if (id_bypass_src_0_0) begin
        ex_reg_rs_lsb_0 <= 2'h0;
      end else if (id_bypass_src_0_1) begin
        ex_reg_rs_lsb_0 <= 2'h1;
      end else if (id_bypass_src_0_2) begin
        ex_reg_rs_lsb_0 <= 2'h2;
      end else begin
        ex_reg_rs_lsb_0 <= 2'h3;
      end
    end
    if (metaReset) begin
      ex_reg_rs_lsb_1 <= 2'h0;
    end else if (~ctrl_killd) begin
      if (_T_1140) begin
        ex_reg_rs_lsb_1 <= id_rs_1[1:0];
      end else if (id_bypass_src_1_0) begin
        ex_reg_rs_lsb_1 <= 2'h0;
      end else if (id_bypass_src_1_1) begin
        ex_reg_rs_lsb_1 <= 2'h1;
      end else if (id_bypass_src_1_2) begin
        ex_reg_rs_lsb_1 <= 2'h2;
      end else begin
        ex_reg_rs_lsb_1 <= 2'h3;
      end
    end
    if (metaReset) begin
      ex_reg_rs_msb_0 <= 62'h0;
    end else if (~ctrl_killd) begin
      if (id_illegal_insn) begin
        ex_reg_rs_msb_0 <= {{32'd0}, inst[31:2]};
      end else if (_T_1132) begin
        ex_reg_rs_msb_0 <= id_rs_0[63:2];
      end
    end
    if (metaReset) begin
      ex_reg_rs_msb_1 <= 62'h0;
    end else if (~ctrl_killd) begin
      if (_T_1140) begin
        ex_reg_rs_msb_1 <= id_rs_1[63:2];
      end
    end
    if (metaReset) begin
      _T_1574 <= 32'h0;
    end else if (reset) begin
      _T_1574 <= 32'h0;
    end else if (_T_1608) begin
      _T_1574 <= _T_1607;
    end else if (ll_wen) begin
      _T_1574 <= _T_1580;
    end
    if (metaReset) begin
      _T_1687 <= 32'h0;
    end else if (reset) begin
      _T_1687 <= 32'h0;
    end else if (_T_1705) begin
      _T_1687 <= _T_1704;
    end else if (_T_1700) begin
      _T_1687 <= _T_1699;
    end else if (_T_1690) begin
      _T_1687 <= _T_1693;
    end
    if (metaReset) begin
      blocked <= 1'h0;
    end else begin
      blocked <= _T_1723 & _T_1725;
    end
    if (metaReset) begin
      _T_1445 <= 1'h0;
    end else begin
      _T_1445 <= div_io_req_ready & div_io_req_valid;
    end
    if (metaReset) begin
      _T_1866 <= 64'h0;
    end else if (ex_reg_rs_bypass_0) begin
      if (_T_1014) begin
        _T_1866 <= io_dmem_resp_bits_data_word_bypass;
      end else if (_T_1012) begin
        _T_1866 <= wb_reg_wdata;
      end else if (_T_1010) begin
        _T_1866 <= mem_reg_wdata;
      end else begin
        _T_1866 <= 64'h0;
      end
    end else begin
      _T_1866 <= _T_1016;
    end
    if (metaReset) begin
      coreMonitorBundle_rd0val <= 64'h0;
    end else begin
      coreMonitorBundle_rd0val <= _T_1866;
    end
    if (metaReset) begin
      _T_1869 <= 64'h0;
    end else if (ex_reg_rs_bypass_1) begin
      if (_T_1021) begin
        _T_1869 <= io_dmem_resp_bits_data_word_bypass;
      end else if (_T_1019) begin
        _T_1869 <= wb_reg_wdata;
      end else if (_T_1017) begin
        _T_1869 <= mem_reg_wdata;
      end else begin
        _T_1869 <= 64'h0;
      end
    end else begin
      _T_1869 <= _T_1023;
    end
    if (metaReset) begin
      coreMonitorBundle_rd1val <= 64'h0;
    end else begin
      coreMonitorBundle_rd1val <= _T_1869;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1849 & ~reset) begin
          $fwrite(32'h80000002,"C%d: %d fetch pc=[%x] inst=[%x] DASM(%x)\n",io_hartid,csr_io_time[31:0],ibuf_io_pc,ibuf_io_inst_0_bits_raw,ibuf_io_inst_0_bits_raw); // @[RocketCore.scala 872:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (csr_io_trace_0_valid & ~reset) begin
          $fwrite(32'h80000002,"C%d: %d [%d] pc=[%x] W[r%d=%x][%d] R[r%d=%x] R[r%d=%x] inst=[%x] DASM(%x)\n",io_hartid,csr_io_time[31:0],coreMonitorBundle_valid,coreMonitorBundle_pc,_T_1872,_T_1873,coreMonitorBundle_wrenx,_T_1875,_T_1877,_T_1879,_T_1881,coreMonitorBundle_inst,coreMonitorBundle_inst); // @[RocketCore.scala 930:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    Rocket_state <= Rocket_xor0;
    if (!(Rocket_cov_read_data)) begin
      Rocket_covSum <= Rocket_covSum + 1'h1;
    end
    if (metaReset) begin
      Rocket_metaAssert <= 1'h0;
    end else begin
      Rocket_metaAssert <= Rocket_metaAssert | Rocket_or0;
    end
  end
  always @(posedge clock) begin
    if(Rocket_cov_write_en & Rocket_cov_write_mask) begin
      Rocket_cov[Rocket_cov_write_addr] <= Rocket_cov_write_data; // @[Coverage map for Rocket]
    end
  end
endmodule
module TLMonitor_35(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [3:0]  io_in_a_bits_size,
  input         io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [7:0]  io_in_a_bits_mask,
  input         io_in_b_ready,
  input         io_in_b_valid,
  input  [2:0]  io_in_b_bits_opcode,
  input  [1:0]  io_in_b_bits_param,
  input  [3:0]  io_in_b_bits_size,
  input         io_in_b_bits_source,
  input  [31:0] io_in_b_bits_address,
  input  [7:0]  io_in_b_bits_mask,
  input         io_in_b_bits_corrupt,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [3:0]  io_in_c_bits_size,
  input         io_in_c_bits_source,
  input  [31:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [3:0]  io_in_d_bits_size,
  input         io_in_d_bits_source,
  input  [1:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_ready,
  input         io_in_e_valid,
  input  [1:0]  io_in_e_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire  _T_7; // @[Parameters.scala 1016:46]
  wire [26:0] _T_9; // @[package.scala 212:77]
  wire [31:0] _GEN_71; // @[Edges.scala 22:16]
  wire [31:0] _T_12; // @[Edges.scala 22:16]
  wire  _T_13; // @[Edges.scala 22:24]
  wire [3:0] _T_16; // @[OneHot.scala 65:12]
  wire [2:0] _T_18; // @[Misc.scala 201:81]
  wire  _T_19; // @[Misc.scala 205:21]
  wire  _T_24; // @[Misc.scala 214:38]
  wire  _T_25; // @[Misc.scala 214:29]
  wire  _T_27; // @[Misc.scala 214:38]
  wire  _T_28; // @[Misc.scala 214:29]
  wire  _T_32; // @[Misc.scala 213:27]
  wire  _T_33; // @[Misc.scala 214:38]
  wire  _T_34; // @[Misc.scala 214:29]
  wire  _T_35; // @[Misc.scala 213:27]
  wire  _T_36; // @[Misc.scala 214:38]
  wire  _T_37; // @[Misc.scala 214:29]
  wire  _T_38; // @[Misc.scala 213:27]
  wire  _T_39; // @[Misc.scala 214:38]
  wire  _T_40; // @[Misc.scala 214:29]
  wire  _T_41; // @[Misc.scala 213:27]
  wire  _T_42; // @[Misc.scala 214:38]
  wire  _T_43; // @[Misc.scala 214:29]
  wire  _T_47; // @[Misc.scala 213:27]
  wire  _T_48; // @[Misc.scala 214:38]
  wire  _T_49; // @[Misc.scala 214:29]
  wire  _T_50; // @[Misc.scala 213:27]
  wire  _T_51; // @[Misc.scala 214:38]
  wire  _T_52; // @[Misc.scala 214:29]
  wire  _T_53; // @[Misc.scala 213:27]
  wire  _T_54; // @[Misc.scala 214:38]
  wire  _T_55; // @[Misc.scala 214:29]
  wire  _T_56; // @[Misc.scala 213:27]
  wire  _T_57; // @[Misc.scala 214:38]
  wire  _T_58; // @[Misc.scala 214:29]
  wire  _T_59; // @[Misc.scala 213:27]
  wire  _T_60; // @[Misc.scala 214:38]
  wire  _T_61; // @[Misc.scala 214:29]
  wire  _T_62; // @[Misc.scala 213:27]
  wire  _T_63; // @[Misc.scala 214:38]
  wire  _T_64; // @[Misc.scala 214:29]
  wire  _T_65; // @[Misc.scala 213:27]
  wire  _T_66; // @[Misc.scala 214:38]
  wire  _T_67; // @[Misc.scala 214:29]
  wire  _T_68; // @[Misc.scala 213:27]
  wire  _T_69; // @[Misc.scala 214:38]
  wire  _T_70; // @[Misc.scala 214:29]
  wire [7:0] _T_77; // @[Cat.scala 29:58]
  wire [32:0] _T_81; // @[Parameters.scala 137:49]
  wire  _T_98; // @[Monitor.scala 82:25]
  wire  _T_100; // @[Parameters.scala 93:42]
  wire  _T_105; // @[Parameters.scala 1066:30]
  wire  _T_115; // @[Parameters.scala 93:42]
  wire [31:0] _T_118; // @[Parameters.scala 137:31]
  wire [32:0] _T_119; // @[Parameters.scala 137:49]
  wire [32:0] _T_121; // @[Parameters.scala 137:52]
  wire  _T_122; // @[Parameters.scala 137:67]
  wire  _T_123; // @[Parameters.scala 601:56]
  wire  _T_126; // @[Parameters.scala 1240:195]
  wire  _T_128; // @[Monitor.scala 44:11]
  wire  _T_133; // @[Parameters.scala 92:48]
  wire  _T_134; // @[Mux.scala 27:72]
  wire  _T_149; // @[Parameters.scala 1255:195]
  wire  _T_151; // @[Monitor.scala 44:11]
  wire  _T_154; // @[Monitor.scala 44:11]
  wire  _T_158; // @[Monitor.scala 44:11]
  wire  _T_161; // @[Monitor.scala 44:11]
  wire  _T_163; // @[Bundles.scala 110:27]
  wire  _T_165; // @[Monitor.scala 44:11]
  wire  _T_168; // @[Monitor.scala 89:31]
  wire  _T_170; // @[Monitor.scala 44:11]
  wire  _T_176; // @[Monitor.scala 93:25]
  wire  _T_245; // @[Monitor.scala 100:31]
  wire  _T_247; // @[Monitor.scala 44:11]
  wire  _T_258; // @[Monitor.scala 105:25]
  wire [31:0] _T_271; // @[Parameters.scala 137:31]
  wire [32:0] _T_272; // @[Parameters.scala 137:49]
  wire [32:0] _T_274; // @[Parameters.scala 137:52]
  wire  _T_275; // @[Parameters.scala 137:67]
  wire  _T_276; // @[Parameters.scala 601:56]
  wire [32:0] _T_284; // @[Parameters.scala 137:52]
  wire  _T_285; // @[Parameters.scala 137:67]
  wire [31:0] _T_286; // @[Parameters.scala 137:31]
  wire [32:0] _T_287; // @[Parameters.scala 137:49]
  wire [32:0] _T_289; // @[Parameters.scala 137:52]
  wire  _T_290; // @[Parameters.scala 137:67]
  wire [31:0] _T_291; // @[Parameters.scala 137:31]
  wire [32:0] _T_292; // @[Parameters.scala 137:49]
  wire [32:0] _T_294; // @[Parameters.scala 137:52]
  wire  _T_295; // @[Parameters.scala 137:67]
  wire [31:0] _T_296; // @[Parameters.scala 137:31]
  wire [32:0] _T_297; // @[Parameters.scala 137:49]
  wire [32:0] _T_299; // @[Parameters.scala 137:52]
  wire  _T_300; // @[Parameters.scala 137:67]
  wire [31:0] _T_301; // @[Parameters.scala 137:31]
  wire [32:0] _T_302; // @[Parameters.scala 137:49]
  wire [32:0] _T_304; // @[Parameters.scala 137:52]
  wire  _T_305; // @[Parameters.scala 137:67]
  wire [32:0] _T_309; // @[Parameters.scala 137:52]
  wire  _T_310; // @[Parameters.scala 137:67]
  wire  _T_311; // @[Parameters.scala 602:42]
  wire  _T_312; // @[Parameters.scala 602:42]
  wire  _T_313; // @[Parameters.scala 602:42]
  wire  _T_314; // @[Parameters.scala 602:42]
  wire  _T_315; // @[Parameters.scala 602:42]
  wire  _T_316; // @[Parameters.scala 601:56]
  wire  _T_318; // @[Parameters.scala 603:30]
  wire  _T_319; // @[Parameters.scala 1243:195]
  wire  _T_321; // @[Monitor.scala 44:11]
  wire  _T_329; // @[Monitor.scala 109:31]
  wire  _T_331; // @[Monitor.scala 44:11]
  wire  _T_333; // @[Monitor.scala 110:30]
  wire  _T_335; // @[Monitor.scala 44:11]
  wire  _T_341; // @[Monitor.scala 114:25]
  wire  _T_384; // @[Parameters.scala 602:42]
  wire  _T_385; // @[Parameters.scala 602:42]
  wire  _T_386; // @[Parameters.scala 602:42]
  wire  _T_387; // @[Parameters.scala 601:56]
  wire  _T_396; // @[Parameters.scala 93:42]
  wire  _T_404; // @[Parameters.scala 601:56]
  wire  _T_406; // @[Parameters.scala 603:30]
  wire  _T_408; // @[Parameters.scala 603:30]
  wire  _T_409; // @[Parameters.scala 1244:195]
  wire  _T_411; // @[Monitor.scala 44:11]
  wire  _T_427; // @[Monitor.scala 122:25]
  wire [7:0] _T_510; // @[Monitor.scala 127:31]
  wire  _T_511; // @[Monitor.scala 127:40]
  wire  _T_513; // @[Monitor.scala 44:11]
  wire  _T_515; // @[Monitor.scala 130:25]
  wire  _T_525; // @[Parameters.scala 93:42]
  wire [32:0] _T_531; // @[Parameters.scala 137:52]
  wire  _T_532; // @[Parameters.scala 137:67]
  wire  _T_538; // @[Parameters.scala 602:42]
  wire  _T_539; // @[Parameters.scala 601:56]
  wire  _T_561; // @[Parameters.scala 1241:195]
  wire  _T_563; // @[Monitor.scala 44:11]
  wire  _T_571; // @[Bundles.scala 140:33]
  wire  _T_573; // @[Monitor.scala 44:11]
  wire  _T_579; // @[Monitor.scala 138:25]
  wire  _T_635; // @[Bundles.scala 147:30]
  wire  _T_637; // @[Monitor.scala 44:11]
  wire  _T_643; // @[Monitor.scala 146:25]
  wire  _T_701; // @[Parameters.scala 1246:195]
  wire  _T_703; // @[Monitor.scala 44:11]
  wire  _T_711; // @[Bundles.scala 160:28]
  wire  _T_713; // @[Monitor.scala 44:11]
  wire  _T_723; // @[Bundles.scala 44:24]
  wire  _T_725; // @[Monitor.scala 51:11]
  wire  _T_730; // @[Parameters.scala 1016:46]
  wire  _T_732; // @[Monitor.scala 310:25]
  wire  _T_734; // @[Monitor.scala 51:11]
  wire  _T_736; // @[Monitor.scala 312:27]
  wire  _T_738; // @[Monitor.scala 51:11]
  wire  _T_740; // @[Monitor.scala 313:28]
  wire  _T_742; // @[Monitor.scala 51:11]
  wire  _T_746; // @[Monitor.scala 51:11]
  wire  _T_750; // @[Monitor.scala 51:11]
  wire  _T_752; // @[Monitor.scala 318:25]
  wire  _T_763; // @[Bundles.scala 104:26]
  wire  _T_765; // @[Monitor.scala 51:11]
  wire  _T_767; // @[Monitor.scala 323:28]
  wire  _T_769; // @[Monitor.scala 51:11]
  wire  _T_780; // @[Monitor.scala 328:25]
  wire  _T_800; // @[Monitor.scala 334:30]
  wire  _T_802; // @[Monitor.scala 51:11]
  wire  _T_809; // @[Monitor.scala 338:25]
  wire  _T_826; // @[Monitor.scala 346:25]
  wire  _T_844; // @[Monitor.scala 354:25]
  wire  _T_861; // @[Bundles.scala 42:24]
  wire  _T_863; // @[Monitor.scala 44:11]
  wire [32:0] _T_868; // @[Parameters.scala 137:49]
  wire [31:0] _T_885; // @[Parameters.scala 137:31]
  wire [32:0] _T_886; // @[Parameters.scala 137:49]
  wire [32:0] _T_888; // @[Parameters.scala 137:52]
  wire  _T_889; // @[Parameters.scala 137:67]
  wire [31:0] _T_890; // @[Parameters.scala 137:31]
  wire [32:0] _T_891; // @[Parameters.scala 137:49]
  wire [32:0] _T_893; // @[Parameters.scala 137:52]
  wire  _T_894; // @[Parameters.scala 137:67]
  wire [31:0] _T_895; // @[Parameters.scala 137:31]
  wire [32:0] _T_896; // @[Parameters.scala 137:49]
  wire [32:0] _T_898; // @[Parameters.scala 137:52]
  wire  _T_899; // @[Parameters.scala 137:67]
  wire [32:0] _T_903; // @[Parameters.scala 137:52]
  wire  _T_904; // @[Parameters.scala 137:67]
  wire [31:0] _T_905; // @[Parameters.scala 137:31]
  wire [32:0] _T_906; // @[Parameters.scala 137:49]
  wire [32:0] _T_908; // @[Parameters.scala 137:52]
  wire  _T_909; // @[Parameters.scala 137:67]
  wire [31:0] _T_910; // @[Parameters.scala 137:31]
  wire [32:0] _T_911; // @[Parameters.scala 137:49]
  wire [32:0] _T_913; // @[Parameters.scala 137:52]
  wire  _T_914; // @[Parameters.scala 137:67]
  wire [31:0] _T_915; // @[Parameters.scala 137:31]
  wire [32:0] _T_916; // @[Parameters.scala 137:49]
  wire [32:0] _T_918; // @[Parameters.scala 137:52]
  wire  _T_919; // @[Parameters.scala 137:67]
  wire  _T_921; // @[Parameters.scala 556:64]
  wire  _T_922; // @[Parameters.scala 556:64]
  wire  _T_923; // @[Parameters.scala 556:64]
  wire  _T_924; // @[Parameters.scala 556:64]
  wire  _T_925; // @[Parameters.scala 556:64]
  wire  _T_926; // @[Parameters.scala 556:64]
  wire [26:0] _T_928; // @[package.scala 212:77]
  wire [31:0] _GEN_72; // @[Edges.scala 22:16]
  wire [31:0] _T_931; // @[Edges.scala 22:16]
  wire  _T_932; // @[Edges.scala 22:24]
  wire [3:0] _T_935; // @[OneHot.scala 65:12]
  wire [2:0] _T_937; // @[Misc.scala 201:81]
  wire  _T_938; // @[Misc.scala 205:21]
  wire  _T_943; // @[Misc.scala 214:38]
  wire  _T_944; // @[Misc.scala 214:29]
  wire  _T_946; // @[Misc.scala 214:38]
  wire  _T_947; // @[Misc.scala 214:29]
  wire  _T_951; // @[Misc.scala 213:27]
  wire  _T_952; // @[Misc.scala 214:38]
  wire  _T_953; // @[Misc.scala 214:29]
  wire  _T_954; // @[Misc.scala 213:27]
  wire  _T_955; // @[Misc.scala 214:38]
  wire  _T_956; // @[Misc.scala 214:29]
  wire  _T_957; // @[Misc.scala 213:27]
  wire  _T_958; // @[Misc.scala 214:38]
  wire  _T_959; // @[Misc.scala 214:29]
  wire  _T_960; // @[Misc.scala 213:27]
  wire  _T_961; // @[Misc.scala 214:38]
  wire  _T_962; // @[Misc.scala 214:29]
  wire  _T_966; // @[Misc.scala 213:27]
  wire  _T_967; // @[Misc.scala 214:38]
  wire  _T_968; // @[Misc.scala 214:29]
  wire  _T_969; // @[Misc.scala 213:27]
  wire  _T_970; // @[Misc.scala 214:38]
  wire  _T_971; // @[Misc.scala 214:29]
  wire  _T_972; // @[Misc.scala 213:27]
  wire  _T_973; // @[Misc.scala 214:38]
  wire  _T_974; // @[Misc.scala 214:29]
  wire  _T_975; // @[Misc.scala 213:27]
  wire  _T_976; // @[Misc.scala 214:38]
  wire  _T_977; // @[Misc.scala 214:29]
  wire  _T_978; // @[Misc.scala 213:27]
  wire  _T_979; // @[Misc.scala 214:38]
  wire  _T_980; // @[Misc.scala 214:29]
  wire  _T_981; // @[Misc.scala 213:27]
  wire  _T_982; // @[Misc.scala 214:38]
  wire  _T_983; // @[Misc.scala 214:29]
  wire  _T_984; // @[Misc.scala 213:27]
  wire  _T_985; // @[Misc.scala 214:38]
  wire  _T_986; // @[Misc.scala 214:29]
  wire  _T_987; // @[Misc.scala 213:27]
  wire  _T_988; // @[Misc.scala 214:38]
  wire  _T_989; // @[Misc.scala 214:29]
  wire [7:0] _T_996; // @[Cat.scala 29:58]
  wire  _T_1004; // @[Monitor.scala 165:113]
  wire  _T_1005; // @[Monitor.scala 167:25]
  wire  _T_1009; // @[Parameters.scala 92:48]
  wire  _T_1010; // @[Mux.scala 27:72]
  wire  _T_1015; // @[Parameters.scala 93:42]
  wire  _T_1025; // @[Parameters.scala 1255:195]
  wire  _T_1027; // @[Monitor.scala 44:11]
  wire  _T_1030; // @[Monitor.scala 44:11]
  wire  _T_1033; // @[Monitor.scala 44:11]
  wire  _T_1036; // @[Monitor.scala 44:11]
  wire  _T_1038; // @[Bundles.scala 104:26]
  wire  _T_1040; // @[Monitor.scala 44:11]
  wire  _T_1042; // @[Monitor.scala 173:30]
  wire  _T_1044; // @[Monitor.scala 44:11]
  wire  _T_1048; // @[Monitor.scala 44:11]
  wire  _T_1050; // @[Monitor.scala 177:25]
  wire  _T_1075; // @[Monitor.scala 182:31]
  wire  _T_1077; // @[Monitor.scala 44:11]
  wire  _T_1087; // @[Monitor.scala 187:25]
  wire  _T_1120; // @[Monitor.scala 196:25]
  wire [7:0] _T_1150; // @[Monitor.scala 202:31]
  wire  _T_1151; // @[Monitor.scala 202:40]
  wire  _T_1153; // @[Monitor.scala 44:11]
  wire  _T_1155; // @[Monitor.scala 205:25]
  wire  _T_1188; // @[Monitor.scala 214:25]
  wire  _T_1221; // @[Monitor.scala 223:25]
  wire  _T_1261; // @[Parameters.scala 1016:46]
  wire [26:0] _T_1263; // @[package.scala 212:77]
  wire [31:0] _GEN_73; // @[Edges.scala 22:16]
  wire [31:0] _T_1266; // @[Edges.scala 22:16]
  wire  _T_1267; // @[Edges.scala 22:24]
  wire [31:0] _T_1268; // @[Parameters.scala 137:31]
  wire [32:0] _T_1269; // @[Parameters.scala 137:49]
  wire [32:0] _T_1271; // @[Parameters.scala 137:52]
  wire  _T_1272; // @[Parameters.scala 137:67]
  wire [31:0] _T_1273; // @[Parameters.scala 137:31]
  wire [32:0] _T_1274; // @[Parameters.scala 137:49]
  wire [32:0] _T_1276; // @[Parameters.scala 137:52]
  wire  _T_1277; // @[Parameters.scala 137:67]
  wire [31:0] _T_1278; // @[Parameters.scala 137:31]
  wire [32:0] _T_1279; // @[Parameters.scala 137:49]
  wire [32:0] _T_1281; // @[Parameters.scala 137:52]
  wire  _T_1282; // @[Parameters.scala 137:67]
  wire [32:0] _T_1284; // @[Parameters.scala 137:49]
  wire [32:0] _T_1286; // @[Parameters.scala 137:52]
  wire  _T_1287; // @[Parameters.scala 137:67]
  wire [31:0] _T_1288; // @[Parameters.scala 137:31]
  wire [32:0] _T_1289; // @[Parameters.scala 137:49]
  wire [32:0] _T_1291; // @[Parameters.scala 137:52]
  wire  _T_1292; // @[Parameters.scala 137:67]
  wire [31:0] _T_1293; // @[Parameters.scala 137:31]
  wire [32:0] _T_1294; // @[Parameters.scala 137:49]
  wire [32:0] _T_1296; // @[Parameters.scala 137:52]
  wire  _T_1297; // @[Parameters.scala 137:67]
  wire [31:0] _T_1298; // @[Parameters.scala 137:31]
  wire [32:0] _T_1299; // @[Parameters.scala 137:49]
  wire [32:0] _T_1301; // @[Parameters.scala 137:52]
  wire  _T_1302; // @[Parameters.scala 137:67]
  wire  _T_1304; // @[Parameters.scala 556:64]
  wire  _T_1305; // @[Parameters.scala 556:64]
  wire  _T_1306; // @[Parameters.scala 556:64]
  wire  _T_1307; // @[Parameters.scala 556:64]
  wire  _T_1308; // @[Parameters.scala 556:64]
  wire  _T_1309; // @[Parameters.scala 556:64]
  wire  _T_1330; // @[Monitor.scala 242:25]
  wire  _T_1332; // @[Monitor.scala 44:11]
  wire  _T_1335; // @[Monitor.scala 44:11]
  wire  _T_1337; // @[Monitor.scala 245:30]
  wire  _T_1339; // @[Monitor.scala 44:11]
  wire  _T_1342; // @[Monitor.scala 44:11]
  wire  _T_1344; // @[Bundles.scala 122:29]
  wire  _T_1346; // @[Monitor.scala 44:11]
  wire  _T_1352; // @[Monitor.scala 251:25]
  wire  _T_1370; // @[Monitor.scala 259:25]
  wire  _T_1372; // @[Parameters.scala 93:42]
  wire  _T_1377; // @[Parameters.scala 1066:30]
  wire  _T_1387; // @[Parameters.scala 93:42]
  wire [32:0] _T_1393; // @[Parameters.scala 137:52]
  wire  _T_1394; // @[Parameters.scala 137:67]
  wire  _T_1395; // @[Parameters.scala 601:56]
  wire  _T_1398; // @[Parameters.scala 1240:195]
  wire  _T_1400; // @[Monitor.scala 44:11]
  wire  _T_1405; // @[Parameters.scala 92:48]
  wire  _T_1406; // @[Mux.scala 27:72]
  wire  _T_1421; // @[Parameters.scala 1255:195]
  wire  _T_1423; // @[Monitor.scala 44:11]
  wire  _T_1435; // @[Bundles.scala 116:29]
  wire  _T_1437; // @[Monitor.scala 44:11]
  wire  _T_1443; // @[Monitor.scala 269:25]
  wire  _T_1512; // @[Monitor.scala 278:25]
  wire  _T_1522; // @[Monitor.scala 282:31]
  wire  _T_1524; // @[Monitor.scala 44:11]
  wire  _T_1530; // @[Monitor.scala 286:25]
  wire  _T_1544; // @[Monitor.scala 293:25]
  wire  _T_1566; // @[Decoupled.scala 40:37]
  wire [8:0] _T_1571; // @[Edges.scala 221:59]
  reg [8:0] _T_1575; // @[Edges.scala 230:27]
  reg [31:0] _RAND_0;
  wire [8:0] _T_1577; // @[Edges.scala 231:28]
  wire  _T_1578; // @[Edges.scala 232:25]
  reg [2:0] _T_1586; // @[Monitor.scala 384:22]
  reg [31:0] _RAND_1;
  reg [2:0] _T_1587; // @[Monitor.scala 385:22]
  reg [31:0] _RAND_2;
  reg [3:0] _T_1588; // @[Monitor.scala 386:22]
  reg [31:0] _RAND_3;
  reg  _T_1589; // @[Monitor.scala 387:22]
  reg [31:0] _RAND_4;
  reg [31:0] _T_1590; // @[Monitor.scala 388:22]
  reg [31:0] _RAND_5;
  wire  _T_1592; // @[Monitor.scala 389:19]
  wire  _T_1593; // @[Monitor.scala 390:32]
  wire  _T_1595; // @[Monitor.scala 44:11]
  wire  _T_1597; // @[Monitor.scala 391:32]
  wire  _T_1599; // @[Monitor.scala 44:11]
  wire  _T_1601; // @[Monitor.scala 392:32]
  wire  _T_1603; // @[Monitor.scala 44:11]
  wire  _T_1605; // @[Monitor.scala 393:32]
  wire  _T_1607; // @[Monitor.scala 44:11]
  wire  _T_1609; // @[Monitor.scala 394:32]
  wire  _T_1611; // @[Monitor.scala 44:11]
  wire  _T_1614; // @[Monitor.scala 396:20]
  wire  _T_1615; // @[Decoupled.scala 40:37]
  wire [26:0] _T_1617; // @[package.scala 212:77]
  wire [8:0] _T_1620; // @[Edges.scala 221:59]
  reg [8:0] _T_1623; // @[Edges.scala 230:27]
  reg [31:0] _RAND_6;
  wire [8:0] _T_1625; // @[Edges.scala 231:28]
  wire  _T_1626; // @[Edges.scala 232:25]
  reg [2:0] _T_1634; // @[Monitor.scala 535:22]
  reg [31:0] _RAND_7;
  reg [1:0] _T_1635; // @[Monitor.scala 536:22]
  reg [31:0] _RAND_8;
  reg [3:0] _T_1636; // @[Monitor.scala 537:22]
  reg [31:0] _RAND_9;
  reg  _T_1637; // @[Monitor.scala 538:22]
  reg [31:0] _RAND_10;
  reg [1:0] _T_1638; // @[Monitor.scala 539:22]
  reg [31:0] _RAND_11;
  reg  _T_1639; // @[Monitor.scala 540:22]
  reg [31:0] _RAND_12;
  wire  _T_1641; // @[Monitor.scala 541:19]
  wire  _T_1642; // @[Monitor.scala 542:29]
  wire  _T_1644; // @[Monitor.scala 51:11]
  wire  _T_1646; // @[Monitor.scala 543:29]
  wire  _T_1648; // @[Monitor.scala 51:11]
  wire  _T_1650; // @[Monitor.scala 544:29]
  wire  _T_1652; // @[Monitor.scala 51:11]
  wire  _T_1654; // @[Monitor.scala 545:29]
  wire  _T_1656; // @[Monitor.scala 51:11]
  wire  _T_1658; // @[Monitor.scala 546:29]
  wire  _T_1660; // @[Monitor.scala 51:11]
  wire  _T_1662; // @[Monitor.scala 547:29]
  wire  _T_1664; // @[Monitor.scala 51:11]
  wire  _T_1667; // @[Monitor.scala 549:20]
  wire  _T_1668; // @[Decoupled.scala 40:37]
  reg [8:0] _T_1677; // @[Edges.scala 230:27]
  reg [31:0] _RAND_13;
  wire [8:0] _T_1679; // @[Edges.scala 231:28]
  wire  _T_1680; // @[Edges.scala 232:25]
  reg [2:0] _T_1688; // @[Monitor.scala 407:22]
  reg [31:0] _RAND_14;
  reg [1:0] _T_1689; // @[Monitor.scala 408:22]
  reg [31:0] _RAND_15;
  reg [3:0] _T_1690; // @[Monitor.scala 409:22]
  reg [31:0] _RAND_16;
  reg  _T_1691; // @[Monitor.scala 410:22]
  reg [31:0] _RAND_17;
  reg [31:0] _T_1692; // @[Monitor.scala 411:22]
  reg [31:0] _RAND_18;
  wire  _T_1694; // @[Monitor.scala 412:19]
  wire  _T_1695; // @[Monitor.scala 413:32]
  wire  _T_1697; // @[Monitor.scala 44:11]
  wire  _T_1699; // @[Monitor.scala 414:32]
  wire  _T_1701; // @[Monitor.scala 44:11]
  wire  _T_1703; // @[Monitor.scala 415:32]
  wire  _T_1705; // @[Monitor.scala 44:11]
  wire  _T_1707; // @[Monitor.scala 416:32]
  wire  _T_1709; // @[Monitor.scala 44:11]
  wire  _T_1711; // @[Monitor.scala 417:32]
  wire  _T_1713; // @[Monitor.scala 44:11]
  wire  _T_1716; // @[Monitor.scala 419:20]
  wire  _T_1717; // @[Decoupled.scala 40:37]
  wire [8:0] _T_1722; // @[Edges.scala 221:59]
  reg [8:0] _T_1725; // @[Edges.scala 230:27]
  reg [31:0] _RAND_19;
  wire [8:0] _T_1727; // @[Edges.scala 231:28]
  wire  _T_1728; // @[Edges.scala 232:25]
  reg [2:0] _T_1736; // @[Monitor.scala 512:22]
  reg [31:0] _RAND_20;
  reg [2:0] _T_1737; // @[Monitor.scala 513:22]
  reg [31:0] _RAND_21;
  reg [3:0] _T_1738; // @[Monitor.scala 514:22]
  reg [31:0] _RAND_22;
  reg  _T_1739; // @[Monitor.scala 515:22]
  reg [31:0] _RAND_23;
  reg [31:0] _T_1740; // @[Monitor.scala 516:22]
  reg [31:0] _RAND_24;
  wire  _T_1742; // @[Monitor.scala 517:19]
  wire  _T_1743; // @[Monitor.scala 518:32]
  wire  _T_1745; // @[Monitor.scala 44:11]
  wire  _T_1747; // @[Monitor.scala 519:32]
  wire  _T_1749; // @[Monitor.scala 44:11]
  wire  _T_1751; // @[Monitor.scala 520:32]
  wire  _T_1753; // @[Monitor.scala 44:11]
  wire  _T_1755; // @[Monitor.scala 521:32]
  wire  _T_1757; // @[Monitor.scala 44:11]
  wire  _T_1759; // @[Monitor.scala 522:32]
  wire  _T_1761; // @[Monitor.scala 44:11]
  wire  _T_1764; // @[Monitor.scala 524:20]
  reg [1:0] inflight; // @[Monitor.scala 611:27]
  reg [31:0] _RAND_25;
  reg [7:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [31:0] _RAND_26;
  reg [15:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [31:0] _RAND_27;
  reg [8:0] _T_1774; // @[Edges.scala 230:27]
  reg [31:0] _RAND_28;
  wire [8:0] _T_1776; // @[Edges.scala 231:28]
  wire  a_first; // @[Edges.scala 232:25]
  reg [8:0] _T_1792; // @[Edges.scala 230:27]
  reg [31:0] _RAND_29;
  wire [8:0] _T_1794; // @[Edges.scala 231:28]
  wire  d_first; // @[Edges.scala 232:25]
  wire [2:0] _GEN_74; // @[Monitor.scala 632:69]
  wire [3:0] _T_1802; // @[Monitor.scala 632:69]
  wire [7:0] _T_1803; // @[Monitor.scala 632:44]
  wire [15:0] _T_1807; // @[Monitor.scala 609:57]
  wire [15:0] _GEN_75; // @[Monitor.scala 632:97]
  wire [15:0] _T_1808; // @[Monitor.scala 632:97]
  wire [15:0] _T_1809; // @[Monitor.scala 632:152]
  wire [3:0] _T_1810; // @[Monitor.scala 636:65]
  wire [15:0] _T_1811; // @[Monitor.scala 636:40]
  wire [15:0] _T_1815; // @[Monitor.scala 609:57]
  wire [15:0] _T_1816; // @[Monitor.scala 636:91]
  wire [15:0] _T_1817; // @[Monitor.scala 636:144]
  wire  _T_1821; // @[Monitor.scala 646:27]
  wire [1:0] _T_1823; // @[OneHot.scala 58:35]
  wire [3:0] _T_1824; // @[Monitor.scala 648:53]
  wire [3:0] _T_1825; // @[Monitor.scala 648:61]
  wire [4:0] _T_1826; // @[Monitor.scala 649:49]
  wire [4:0] _T_1827; // @[Monitor.scala 649:57]
  wire [2:0] _GEN_78; // @[Monitor.scala 650:72]
  wire [3:0] _T_1828; // @[Monitor.scala 650:72]
  wire [3:0] a_opcodes_set_interm; // @[Monitor.scala 646:72]
  wire [18:0] _GEN_79; // @[Monitor.scala 650:47]
  wire [18:0] _T_1829; // @[Monitor.scala 650:47]
  wire [3:0] _T_1830; // @[Monitor.scala 651:68]
  wire [4:0] a_sizes_set_interm; // @[Monitor.scala 646:72]
  wire [19:0] _GEN_80; // @[Monitor.scala 651:43]
  wire [19:0] _T_1831; // @[Monitor.scala 651:43]
  wire [1:0] _T_1832; // @[Monitor.scala 652:26]
  wire  _T_1836; // @[Monitor.scala 44:11]
  wire [1:0] a_set; // @[Monitor.scala 646:72]
  wire [18:0] _GEN_30; // @[Monitor.scala 646:72]
  wire [19:0] _GEN_31; // @[Monitor.scala 646:72]
  wire  _T_1840; // @[Monitor.scala 663:27]
  wire  _T_1843; // @[Monitor.scala 663:72]
  wire [1:0] _T_1844; // @[OneHot.scala 58:35]
  wire [30:0] _GEN_82; // @[Monitor.scala 665:76]
  wire [30:0] _T_1850; // @[Monitor.scala 665:76]
  wire [30:0] _GEN_83; // @[Monitor.scala 666:72]
  wire [30:0] _T_1856; // @[Monitor.scala 666:72]
  wire [1:0] d_clr; // @[Monitor.scala 663:91]
  wire [30:0] _GEN_33; // @[Monitor.scala 663:91]
  wire [30:0] _GEN_34; // @[Monitor.scala 663:91]
  wire  _T_1857; // @[Monitor.scala 668:26]
  wire  _T_1860; // @[Monitor.scala 668:71]
  wire [1:0] _T_1861; // @[Monitor.scala 669:25]
  wire  _T_1863; // @[Monitor.scala 669:93]
  wire  _T_1864; // @[Monitor.scala 669:68]
  wire  _T_1865; // @[Monitor.scala 669:142]
  wire  _T_1866; // @[Monitor.scala 669:119]
  wire  _T_1867; // @[Monitor.scala 669:166]
  wire  _T_1868; // @[Monitor.scala 669:49]
  wire  _T_1870; // @[Monitor.scala 51:11]
  wire [3:0] a_opcode_lookup; // @[Monitor.scala 632:21]
  wire [2:0] _GEN_37; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_38; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_39; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_40; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_41; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_42; // @[Monitor.scala 670:37]
  wire  _T_1873; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_49; // @[Monitor.scala 670:96]
  wire [2:0] _GEN_50; // @[Monitor.scala 670:96]
  wire  _T_1875; // @[Monitor.scala 670:96]
  wire  _T_1876; // @[Monitor.scala 670:71]
  wire [2:0] _GEN_53; // @[Monitor.scala 671:60]
  wire [2:0] _GEN_54; // @[Monitor.scala 671:60]
  wire [2:0] _GEN_55; // @[Monitor.scala 671:60]
  wire [2:0] _GEN_56; // @[Monitor.scala 671:60]
  wire [2:0] _GEN_57; // @[Monitor.scala 671:60]
  wire [2:0] _GEN_58; // @[Monitor.scala 671:60]
  wire  _T_1877; // @[Monitor.scala 671:60]
  wire [2:0] _GEN_65; // @[Monitor.scala 671:124]
  wire [2:0] _GEN_66; // @[Monitor.scala 671:124]
  wire  _T_1878; // @[Monitor.scala 671:124]
  wire  _T_1879; // @[Monitor.scala 671:99]
  wire  _T_1880; // @[Monitor.scala 671:34]
  wire  _T_1881; // @[Monitor.scala 671:15]
  wire  _T_1883; // @[Monitor.scala 51:11]
  wire [7:0] a_size_lookup; // @[Monitor.scala 636:19]
  wire [7:0] _GEN_84; // @[Monitor.scala 673:34]
  wire  _T_1885; // @[Monitor.scala 673:34]
  wire  _T_1887; // @[Monitor.scala 673:72]
  wire  _T_1888; // @[Monitor.scala 673:53]
  wire  _T_1890; // @[Monitor.scala 51:11]
  wire  _T_1893; // @[Monitor.scala 675:36]
  wire  _T_1894; // @[Monitor.scala 675:47]
  wire  _T_1896; // @[Monitor.scala 675:65]
  wire  _T_1898; // @[Monitor.scala 675:116]
  wire  _T_1900; // @[Monitor.scala 676:32]
  wire  _T_1902; // @[Monitor.scala 51:11]
  wire  _T_1904; // @[Monitor.scala 680:20]
  wire  _T_1905; // @[Monitor.scala 680:40]
  wire  _T_1907; // @[Monitor.scala 680:30]
  wire  _T_1909; // @[Monitor.scala 51:11]
  wire [1:0] _T_1911; // @[Monitor.scala 683:27]
  wire [1:0] _T_1913; // @[Monitor.scala 683:36]
  wire [7:0] a_opcodes_set; // @[Monitor.scala 650:21]
  wire [7:0] _T_1914; // @[Monitor.scala 684:43]
  wire [7:0] d_opcodes_clr; // @[Monitor.scala 665:21]
  wire [7:0] _T_1916; // @[Monitor.scala 684:60]
  wire [15:0] a_sizes_set; // @[Monitor.scala 651:19]
  wire [15:0] _T_1917; // @[Monitor.scala 685:39]
  wire [15:0] d_sizes_clr; // @[Monitor.scala 666:19]
  wire [15:0] _T_1919; // @[Monitor.scala 685:54]
  reg [3:0] _T_1935; // @[Monitor.scala 697:27]
  reg [31:0] _RAND_30;
  reg [8:0] _T_1944; // @[Edges.scala 230:27]
  reg [31:0] _RAND_31;
  wire [8:0] _T_1946; // @[Edges.scala 231:28]
  wire  _T_1947; // @[Edges.scala 232:25]
  wire  _T_1957; // @[Monitor.scala 703:27]
  wire  _T_1961; // @[Edges.scala 72:40]
  wire  _T_1962; // @[Monitor.scala 703:38]
  wire [3:0] _T_1963; // @[OneHot.scala 58:35]
  wire [3:0] _T_1964; // @[Monitor.scala 705:23]
  wire  _T_1968; // @[Monitor.scala 51:11]
  wire [3:0] _GEN_69; // @[Monitor.scala 703:72]
  wire  _T_1971; // @[Decoupled.scala 40:37]
  wire [3:0] _T_1974; // @[OneHot.scala 58:35]
  wire [3:0] _T_1975; // @[Monitor.scala 711:24]
  wire [3:0] _T_1976; // @[Monitor.scala 711:35]
  wire  _T_1979; // @[Monitor.scala 44:11]
  wire [3:0] _GEN_70; // @[Monitor.scala 709:73]
  wire [3:0] _T_1981; // @[Monitor.scala 716:27]
  wire [3:0] _T_1983; // @[Monitor.scala 716:36]
  wire  _GEN_85; // @[Monitor.scala 44:11]
  wire  _GEN_99; // @[Monitor.scala 44:11]
  wire  _GEN_115; // @[Monitor.scala 44:11]
  wire  _GEN_125; // @[Monitor.scala 44:11]
  wire  _GEN_135; // @[Monitor.scala 44:11]
  wire  _GEN_145; // @[Monitor.scala 44:11]
  wire  _GEN_155; // @[Monitor.scala 44:11]
  wire  _GEN_165; // @[Monitor.scala 44:11]
  wire  _GEN_175; // @[Monitor.scala 51:11]
  wire  _GEN_185; // @[Monitor.scala 51:11]
  wire  _GEN_195; // @[Monitor.scala 51:11]
  wire  _GEN_205; // @[Monitor.scala 51:11]
  wire  _GEN_211; // @[Monitor.scala 51:11]
  wire  _GEN_217; // @[Monitor.scala 51:11]
  wire  _GEN_223; // @[Monitor.scala 44:11]
  wire  _GEN_237; // @[Monitor.scala 44:11]
  wire  _GEN_251; // @[Monitor.scala 44:11]
  wire  _GEN_263; // @[Monitor.scala 44:11]
  wire  _GEN_275; // @[Monitor.scala 44:11]
  wire  _GEN_285; // @[Monitor.scala 44:11]
  wire  _GEN_295; // @[Monitor.scala 44:11]
  wire  _GEN_307; // @[Monitor.scala 44:11]
  wire  _GEN_317; // @[Monitor.scala 44:11]
  wire  _GEN_327; // @[Monitor.scala 44:11]
  wire  _GEN_339; // @[Monitor.scala 44:11]
  wire  _GEN_351; // @[Monitor.scala 44:11]
  wire  _GEN_359; // @[Monitor.scala 44:11]
  wire  _GEN_367; // @[Monitor.scala 44:11]
  wire [29:0] TLMonitor_35_covSum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  stopEn4;
  wire  stopEn5;
  wire  stopEn6;
  wire  stopEn7;
  wire  stopEn8;
  wire  stopEn9;
  wire  stopEn10;
  wire  stopEn11;
  wire  stopEn12;
  wire  stopEn13;
  wire  stopEn14;
  wire  stopEn15;
  wire  stopEn16;
  wire  stopEn17;
  wire  stopEn18;
  wire  stopEn19;
  wire  stopEn20;
  wire  stopEn21;
  wire  stopEn22;
  wire  stopEn23;
  wire  stopEn24;
  wire  stopEn25;
  wire  stopEn26;
  wire  stopEn27;
  wire  stopEn28;
  wire  stopEn29;
  wire  stopEn30;
  wire  stopEn31;
  wire  stopEn32;
  wire  stopEn33;
  wire  stopEn34;
  wire  stopEn35;
  wire  stopEn36;
  wire  stopEn37;
  wire  stopEn38;
  wire  stopEn39;
  wire  stopEn40;
  wire  stopEn41;
  wire  stopEn42;
  wire  stopEn43;
  wire  stopEn44;
  wire  stopEn45;
  wire  stopEn46;
  wire  stopEn47;
  wire  stopEn48;
  wire  stopEn49;
  wire  stopEn50;
  wire  stopEn51;
  wire  stopEn52;
  wire  stopEn53;
  wire  stopEn54;
  wire  stopEn55;
  wire  stopEn56;
  wire  stopEn57;
  wire  stopEn58;
  wire  stopEn59;
  wire  stopEn60;
  wire  stopEn61;
  wire  stopEn62;
  wire  stopEn63;
  wire  stopEn64;
  wire  stopEn65;
  wire  stopEn66;
  wire  stopEn67;
  wire  stopEn68;
  wire  stopEn69;
  wire  stopEn70;
  wire  stopEn71;
  wire  stopEn72;
  wire  stopEn73;
  wire  stopEn74;
  wire  stopEn75;
  wire  stopEn76;
  wire  stopEn77;
  wire  stopEn78;
  wire  stopEn79;
  wire  stopEn80;
  wire  stopEn81;
  wire  stopEn82;
  wire  stopEn83;
  wire  stopEn84;
  wire  stopEn85;
  wire  stopEn86;
  wire  stopEn87;
  wire  stopEn88;
  wire  stopEn89;
  wire  stopEn90;
  wire  stopEn91;
  wire  stopEn92;
  wire  stopEn93;
  wire  stopEn94;
  wire  stopEn95;
  wire  stopEn96;
  wire  stopEn97;
  wire  stopEn98;
  wire  stopEn99;
  wire  stopEn100;
  wire  stopEn101;
  wire  stopEn102;
  wire  stopEn103;
  wire  stopEn104;
  wire  stopEn105;
  wire  stopEn106;
  wire  stopEn107;
  wire  stopEn108;
  wire  stopEn109;
  wire  stopEn110;
  wire  stopEn111;
  wire  stopEn112;
  wire  stopEn113;
  wire  stopEn114;
  wire  stopEn115;
  wire  stopEn116;
  wire  stopEn117;
  wire  stopEn118;
  wire  stopEn119;
  wire  stopEn120;
  wire  stopEn121;
  wire  stopEn122;
  wire  stopEn123;
  wire  stopEn124;
  wire  stopEn125;
  wire  stopEn126;
  wire  stopEn127;
  wire  stopEn128;
  wire  stopEn129;
  wire  stopEn130;
  wire  stopEn131;
  wire  stopEn132;
  wire  stopEn133;
  wire  stopEn134;
  wire  stopEn135;
  wire  stopEn136;
  wire  stopEn137;
  wire  stopEn138;
  wire  stopEn139;
  wire  stopEn140;
  wire  stopEn141;
  wire  stopEn142;
  wire  stopEn143;
  wire  stopEn144;
  wire  stopEn145;
  wire  stopEn146;
  wire  stopEn147;
  wire  stopEn148;
  wire  stopEn149;
  wire  stopEn150;
  wire  stopEn151;
  wire  stopEn152;
  wire  stopEn153;
  wire  stopEn154;
  wire  stopEn155;
  wire  stopEn156;
  wire  stopEn157;
  wire  stopEn158;
  wire  stopEn159;
  wire  stopEn160;
  wire  stopEn161;
  wire  stopEn162;
  wire  stopEn163;
  wire  stopEn164;
  wire  stopEn165;
  wire  stopEn166;
  wire  stopEn167;
  wire  stopEn168;
  wire  stopEn169;
  wire  stopEn170;
  wire  stopEn171;
  wire  stopEn172;
  wire  stopEn173;
  wire  stopEn174;
  wire  stopEn175;
  wire  TLMonitor_35_or63;
  wire  TLMonitor_35_or130;
  wire  TLMonitor_35_or64;
  wire  TLMonitor_35_or31;
  wire  TLMonitor_35_or132;
  wire  TLMonitor_35_or65;
  wire  TLMonitor_35_or134;
  wire  TLMonitor_35_or66;
  wire  TLMonitor_35_or32;
  wire  TLMonitor_35_or15;
  wire  TLMonitor_35_or67;
  wire  TLMonitor_35_or138;
  wire  TLMonitor_35_or68;
  wire  TLMonitor_35_or33;
  wire  TLMonitor_35_or140;
  wire  TLMonitor_35_or69;
  wire  TLMonitor_35_or142;
  wire  TLMonitor_35_or70;
  wire  TLMonitor_35_or34;
  wire  TLMonitor_35_or16;
  wire  TLMonitor_35_or7;
  wire  TLMonitor_35_or71;
  wire  TLMonitor_35_or146;
  wire  TLMonitor_35_or72;
  wire  TLMonitor_35_or35;
  wire  TLMonitor_35_or148;
  wire  TLMonitor_35_or73;
  wire  TLMonitor_35_or150;
  wire  TLMonitor_35_or74;
  wire  TLMonitor_35_or36;
  wire  TLMonitor_35_or17;
  wire  TLMonitor_35_or75;
  wire  TLMonitor_35_or154;
  wire  TLMonitor_35_or76;
  wire  TLMonitor_35_or37;
  wire  TLMonitor_35_or156;
  wire  TLMonitor_35_or77;
  wire  TLMonitor_35_or158;
  wire  TLMonitor_35_or78;
  wire  TLMonitor_35_or38;
  wire  TLMonitor_35_or18;
  wire  TLMonitor_35_or8;
  wire  TLMonitor_35_or3;
  wire  TLMonitor_35_or79;
  wire  TLMonitor_35_or162;
  wire  TLMonitor_35_or80;
  wire  TLMonitor_35_or39;
  wire  TLMonitor_35_or164;
  wire  TLMonitor_35_or81;
  wire  TLMonitor_35_or166;
  wire  TLMonitor_35_or82;
  wire  TLMonitor_35_or40;
  wire  TLMonitor_35_or19;
  wire  TLMonitor_35_or83;
  wire  TLMonitor_35_or170;
  wire  TLMonitor_35_or84;
  wire  TLMonitor_35_or41;
  wire  TLMonitor_35_or172;
  wire  TLMonitor_35_or85;
  wire  TLMonitor_35_or174;
  wire  TLMonitor_35_or86;
  wire  TLMonitor_35_or42;
  wire  TLMonitor_35_or20;
  wire  TLMonitor_35_or9;
  wire  TLMonitor_35_or87;
  wire  TLMonitor_35_or178;
  wire  TLMonitor_35_or88;
  wire  TLMonitor_35_or43;
  wire  TLMonitor_35_or180;
  wire  TLMonitor_35_or89;
  wire  TLMonitor_35_or182;
  wire  TLMonitor_35_or90;
  wire  TLMonitor_35_or44;
  wire  TLMonitor_35_or21;
  wire  TLMonitor_35_or91;
  wire  TLMonitor_35_or186;
  wire  TLMonitor_35_or92;
  wire  TLMonitor_35_or45;
  wire  TLMonitor_35_or188;
  wire  TLMonitor_35_or93;
  wire  TLMonitor_35_or190;
  wire  TLMonitor_35_or94;
  wire  TLMonitor_35_or46;
  wire  TLMonitor_35_or22;
  wire  TLMonitor_35_or10;
  wire  TLMonitor_35_or4;
  wire  TLMonitor_35_or1;
  wire  TLMonitor_35_or95;
  wire  TLMonitor_35_or194;
  wire  TLMonitor_35_or96;
  wire  TLMonitor_35_or47;
  wire  TLMonitor_35_or196;
  wire  TLMonitor_35_or97;
  wire  TLMonitor_35_or198;
  wire  TLMonitor_35_or98;
  wire  TLMonitor_35_or48;
  wire  TLMonitor_35_or23;
  wire  TLMonitor_35_or99;
  wire  TLMonitor_35_or202;
  wire  TLMonitor_35_or100;
  wire  TLMonitor_35_or49;
  wire  TLMonitor_35_or204;
  wire  TLMonitor_35_or101;
  wire  TLMonitor_35_or206;
  wire  TLMonitor_35_or102;
  wire  TLMonitor_35_or50;
  wire  TLMonitor_35_or24;
  wire  TLMonitor_35_or11;
  wire  TLMonitor_35_or103;
  wire  TLMonitor_35_or210;
  wire  TLMonitor_35_or104;
  wire  TLMonitor_35_or51;
  wire  TLMonitor_35_or212;
  wire  TLMonitor_35_or105;
  wire  TLMonitor_35_or214;
  wire  TLMonitor_35_or106;
  wire  TLMonitor_35_or52;
  wire  TLMonitor_35_or25;
  wire  TLMonitor_35_or107;
  wire  TLMonitor_35_or218;
  wire  TLMonitor_35_or108;
  wire  TLMonitor_35_or53;
  wire  TLMonitor_35_or220;
  wire  TLMonitor_35_or109;
  wire  TLMonitor_35_or222;
  wire  TLMonitor_35_or110;
  wire  TLMonitor_35_or54;
  wire  TLMonitor_35_or26;
  wire  TLMonitor_35_or12;
  wire  TLMonitor_35_or5;
  wire  TLMonitor_35_or111;
  wire  TLMonitor_35_or226;
  wire  TLMonitor_35_or112;
  wire  TLMonitor_35_or55;
  wire  TLMonitor_35_or228;
  wire  TLMonitor_35_or113;
  wire  TLMonitor_35_or230;
  wire  TLMonitor_35_or114;
  wire  TLMonitor_35_or56;
  wire  TLMonitor_35_or27;
  wire  TLMonitor_35_or115;
  wire  TLMonitor_35_or234;
  wire  TLMonitor_35_or116;
  wire  TLMonitor_35_or57;
  wire  TLMonitor_35_or236;
  wire  TLMonitor_35_or117;
  wire  TLMonitor_35_or238;
  wire  TLMonitor_35_or118;
  wire  TLMonitor_35_or58;
  wire  TLMonitor_35_or28;
  wire  TLMonitor_35_or13;
  wire  TLMonitor_35_or119;
  wire  TLMonitor_35_or242;
  wire  TLMonitor_35_or120;
  wire  TLMonitor_35_or59;
  wire  TLMonitor_35_or244;
  wire  TLMonitor_35_or121;
  wire  TLMonitor_35_or246;
  wire  TLMonitor_35_or122;
  wire  TLMonitor_35_or60;
  wire  TLMonitor_35_or29;
  wire  TLMonitor_35_or123;
  wire  TLMonitor_35_or250;
  wire  TLMonitor_35_or124;
  wire  TLMonitor_35_or61;
  wire  TLMonitor_35_or252;
  wire  TLMonitor_35_or125;
  wire  TLMonitor_35_or254;
  wire  TLMonitor_35_or126;
  wire  TLMonitor_35_or62;
  wire  TLMonitor_35_or30;
  wire  TLMonitor_35_or14;
  wire  TLMonitor_35_or6;
  wire  TLMonitor_35_or2;
  wire  TLMonitor_35_or0;
  reg  TLMonitor_35_metaAssert;
  reg [31:0] _RAND_32;
  assign _T_7 = ~io_in_a_bits_source | io_in_a_bits_source; // @[Parameters.scala 1016:46]
  assign _T_9 = 27'hfff << io_in_a_bits_size; // @[package.scala 212:77]
  assign _GEN_71 = {{20'd0}, ~_T_9[11:0]}; // @[Edges.scala 22:16]
  assign _T_12 = io_in_a_bits_address & _GEN_71; // @[Edges.scala 22:16]
  assign _T_13 = _T_12 == 32'h0; // @[Edges.scala 22:24]
  assign _T_16 = 4'h1 << io_in_a_bits_size[1:0]; // @[OneHot.scala 65:12]
  assign _T_18 = _T_16[2:0] | 3'h1; // @[Misc.scala 201:81]
  assign _T_19 = io_in_a_bits_size >= 4'h3; // @[Misc.scala 205:21]
  assign _T_24 = _T_18[2] & ~io_in_a_bits_address[2]; // @[Misc.scala 214:38]
  assign _T_25 = _T_19 | _T_24; // @[Misc.scala 214:29]
  assign _T_27 = _T_18[2] & io_in_a_bits_address[2]; // @[Misc.scala 214:38]
  assign _T_28 = _T_19 | _T_27; // @[Misc.scala 214:29]
  assign _T_32 = ~io_in_a_bits_address[2] & ~io_in_a_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_33 = _T_18[1] & _T_32; // @[Misc.scala 214:38]
  assign _T_34 = _T_25 | _T_33; // @[Misc.scala 214:29]
  assign _T_35 = ~io_in_a_bits_address[2] & io_in_a_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_36 = _T_18[1] & _T_35; // @[Misc.scala 214:38]
  assign _T_37 = _T_25 | _T_36; // @[Misc.scala 214:29]
  assign _T_38 = io_in_a_bits_address[2] & ~io_in_a_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_39 = _T_18[1] & _T_38; // @[Misc.scala 214:38]
  assign _T_40 = _T_28 | _T_39; // @[Misc.scala 214:29]
  assign _T_41 = io_in_a_bits_address[2] & io_in_a_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_42 = _T_18[1] & _T_41; // @[Misc.scala 214:38]
  assign _T_43 = _T_28 | _T_42; // @[Misc.scala 214:29]
  assign _T_47 = _T_32 & ~io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_48 = _T_18[0] & _T_47; // @[Misc.scala 214:38]
  assign _T_49 = _T_34 | _T_48; // @[Misc.scala 214:29]
  assign _T_50 = _T_32 & io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_51 = _T_18[0] & _T_50; // @[Misc.scala 214:38]
  assign _T_52 = _T_34 | _T_51; // @[Misc.scala 214:29]
  assign _T_53 = _T_35 & ~io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_54 = _T_18[0] & _T_53; // @[Misc.scala 214:38]
  assign _T_55 = _T_37 | _T_54; // @[Misc.scala 214:29]
  assign _T_56 = _T_35 & io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_57 = _T_18[0] & _T_56; // @[Misc.scala 214:38]
  assign _T_58 = _T_37 | _T_57; // @[Misc.scala 214:29]
  assign _T_59 = _T_38 & ~io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_60 = _T_18[0] & _T_59; // @[Misc.scala 214:38]
  assign _T_61 = _T_40 | _T_60; // @[Misc.scala 214:29]
  assign _T_62 = _T_38 & io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_63 = _T_18[0] & _T_62; // @[Misc.scala 214:38]
  assign _T_64 = _T_40 | _T_63; // @[Misc.scala 214:29]
  assign _T_65 = _T_41 & ~io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_66 = _T_18[0] & _T_65; // @[Misc.scala 214:38]
  assign _T_67 = _T_43 | _T_66; // @[Misc.scala 214:29]
  assign _T_68 = _T_41 & io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_69 = _T_18[0] & _T_68; // @[Misc.scala 214:38]
  assign _T_70 = _T_43 | _T_69; // @[Misc.scala 214:29]
  assign _T_77 = {_T_70,_T_67,_T_64,_T_61,_T_58,_T_55,_T_52,_T_49}; // @[Cat.scala 29:58]
  assign _T_81 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49]
  assign _T_98 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 82:25]
  assign _T_100 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 93:42]
  assign _T_105 = _T_100 & _T_7; // @[Parameters.scala 1066:30]
  assign _T_115 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 93:42]
  assign _T_118 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  assign _T_119 = {1'b0,$signed(_T_118)}; // @[Parameters.scala 137:49]
  assign _T_121 = $signed(_T_119) & 33'sh80000000; // @[Parameters.scala 137:52]
  assign _T_122 = $signed(_T_121) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_123 = _T_115 & _T_122; // @[Parameters.scala 601:56]
  assign _T_126 = _T_105 & _T_123; // @[Parameters.scala 1240:195]
  assign _T_128 = _T_126 | reset; // @[Monitor.scala 44:11]
  assign _T_133 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 92:48]
  assign _T_134 = ~io_in_a_bits_source & _T_133; // @[Mux.scala 27:72]
  assign _T_149 = _T_134 & _T_100; // @[Parameters.scala 1255:195]
  assign _T_151 = _T_149 | reset; // @[Monitor.scala 44:11]
  assign _T_154 = _T_7 | reset; // @[Monitor.scala 44:11]
  assign _T_158 = _T_19 | reset; // @[Monitor.scala 44:11]
  assign _T_161 = _T_13 | reset; // @[Monitor.scala 44:11]
  assign _T_163 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 110:27]
  assign _T_165 = _T_163 | reset; // @[Monitor.scala 44:11]
  assign _T_168 = ~io_in_a_bits_mask == 8'h0; // @[Monitor.scala 89:31]
  assign _T_170 = _T_168 | reset; // @[Monitor.scala 44:11]
  assign _T_176 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 93:25]
  assign _T_245 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 100:31]
  assign _T_247 = _T_245 | reset; // @[Monitor.scala 44:11]
  assign _T_258 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 105:25]
  assign _T_271 = io_in_a_bits_address ^ 32'h2000; // @[Parameters.scala 137:31]
  assign _T_272 = {1'b0,$signed(_T_271)}; // @[Parameters.scala 137:49]
  assign _T_274 = $signed(_T_272) & 33'shca012000; // @[Parameters.scala 137:52]
  assign _T_275 = $signed(_T_274) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_276 = _T_100 & _T_275; // @[Parameters.scala 601:56]
  assign _T_284 = $signed(_T_81) & 33'shca012000; // @[Parameters.scala 137:52]
  assign _T_285 = $signed(_T_284) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_286 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31]
  assign _T_287 = {1'b0,$signed(_T_286)}; // @[Parameters.scala 137:49]
  assign _T_289 = $signed(_T_287) & 33'shca010000; // @[Parameters.scala 137:52]
  assign _T_290 = $signed(_T_289) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_291 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31]
  assign _T_292 = {1'b0,$signed(_T_291)}; // @[Parameters.scala 137:49]
  assign _T_294 = $signed(_T_292) & 33'shca010000; // @[Parameters.scala 137:52]
  assign _T_295 = $signed(_T_294) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_296 = io_in_a_bits_address ^ 32'h8000000; // @[Parameters.scala 137:31]
  assign _T_297 = {1'b0,$signed(_T_296)}; // @[Parameters.scala 137:49]
  assign _T_299 = $signed(_T_297) & 33'shc8000000; // @[Parameters.scala 137:52]
  assign _T_300 = $signed(_T_299) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_301 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  assign _T_302 = {1'b0,$signed(_T_301)}; // @[Parameters.scala 137:49]
  assign _T_304 = $signed(_T_302) & 33'shc0000000; // @[Parameters.scala 137:52]
  assign _T_305 = $signed(_T_304) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_309 = $signed(_T_119) & 33'shc0000000; // @[Parameters.scala 137:52]
  assign _T_310 = $signed(_T_309) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_311 = _T_285 | _T_290; // @[Parameters.scala 602:42]
  assign _T_312 = _T_311 | _T_295; // @[Parameters.scala 602:42]
  assign _T_313 = _T_312 | _T_300; // @[Parameters.scala 602:42]
  assign _T_314 = _T_313 | _T_305; // @[Parameters.scala 602:42]
  assign _T_315 = _T_314 | _T_310; // @[Parameters.scala 602:42]
  assign _T_316 = _T_115 & _T_315; // @[Parameters.scala 601:56]
  assign _T_318 = _T_276 | _T_316; // @[Parameters.scala 603:30]
  assign _T_319 = _T_105 & _T_318; // @[Parameters.scala 1243:195]
  assign _T_321 = _T_319 | reset; // @[Monitor.scala 44:11]
  assign _T_329 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31]
  assign _T_331 = _T_329 | reset; // @[Monitor.scala 44:11]
  assign _T_333 = io_in_a_bits_mask == _T_77; // @[Monitor.scala 110:30]
  assign _T_335 = _T_333 | reset; // @[Monitor.scala 44:11]
  assign _T_341 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  assign _T_384 = _T_285 | _T_295; // @[Parameters.scala 602:42]
  assign _T_385 = _T_384 | _T_300; // @[Parameters.scala 602:42]
  assign _T_386 = _T_385 | _T_310; // @[Parameters.scala 602:42]
  assign _T_387 = _T_115 & _T_386; // @[Parameters.scala 601:56]
  assign _T_396 = io_in_a_bits_size <= 4'h8; // @[Parameters.scala 93:42]
  assign _T_404 = _T_396 & _T_305; // @[Parameters.scala 601:56]
  assign _T_406 = _T_276 | _T_387; // @[Parameters.scala 603:30]
  assign _T_408 = _T_406 | _T_404; // @[Parameters.scala 603:30]
  assign _T_409 = _T_105 & _T_408; // @[Parameters.scala 1244:195]
  assign _T_411 = _T_409 | reset; // @[Monitor.scala 44:11]
  assign _T_427 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  assign _T_510 = io_in_a_bits_mask & ~_T_77; // @[Monitor.scala 127:31]
  assign _T_511 = _T_510 == 8'h0; // @[Monitor.scala 127:40]
  assign _T_513 = _T_511 | reset; // @[Monitor.scala 44:11]
  assign _T_515 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  assign _T_525 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 93:42]
  assign _T_531 = $signed(_T_81) & 33'shc8010000; // @[Parameters.scala 137:52]
  assign _T_532 = $signed(_T_531) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_538 = _T_532 | _T_300; // @[Parameters.scala 602:42]
  assign _T_539 = _T_525 & _T_538; // @[Parameters.scala 601:56]
  assign _T_561 = _T_105 & _T_539; // @[Parameters.scala 1241:195]
  assign _T_563 = _T_561 | reset; // @[Monitor.scala 44:11]
  assign _T_571 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 140:33]
  assign _T_573 = _T_571 | reset; // @[Monitor.scala 44:11]
  assign _T_579 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  assign _T_635 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 147:30]
  assign _T_637 = _T_635 | reset; // @[Monitor.scala 44:11]
  assign _T_643 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  assign _T_701 = _T_105 & _T_276; // @[Parameters.scala 1246:195]
  assign _T_703 = _T_701 | reset; // @[Monitor.scala 44:11]
  assign _T_711 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 160:28]
  assign _T_713 = _T_711 | reset; // @[Monitor.scala 44:11]
  assign _T_723 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 44:24]
  assign _T_725 = _T_723 | reset; // @[Monitor.scala 51:11]
  assign _T_730 = ~io_in_d_bits_source | io_in_d_bits_source; // @[Parameters.scala 1016:46]
  assign _T_732 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  assign _T_734 = _T_730 | reset; // @[Monitor.scala 51:11]
  assign _T_736 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27]
  assign _T_738 = _T_736 | reset; // @[Monitor.scala 51:11]
  assign _T_740 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  assign _T_742 = _T_740 | reset; // @[Monitor.scala 51:11]
  assign _T_746 = ~io_in_d_bits_corrupt | reset; // @[Monitor.scala 51:11]
  assign _T_750 = ~io_in_d_bits_denied | reset; // @[Monitor.scala 51:11]
  assign _T_752 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  assign _T_763 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 104:26]
  assign _T_765 = _T_763 | reset; // @[Monitor.scala 51:11]
  assign _T_767 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  assign _T_769 = _T_767 | reset; // @[Monitor.scala 51:11]
  assign _T_780 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  assign _T_800 = ~io_in_d_bits_denied | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  assign _T_802 = _T_800 | reset; // @[Monitor.scala 51:11]
  assign _T_809 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  assign _T_826 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  assign _T_844 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  assign _T_861 = io_in_b_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  assign _T_863 = _T_861 | reset; // @[Monitor.scala 44:11]
  assign _T_868 = {1'b0,$signed(io_in_b_bits_address)}; // @[Parameters.scala 137:49]
  assign _T_885 = io_in_b_bits_address ^ 32'h3000; // @[Parameters.scala 137:31]
  assign _T_886 = {1'b0,$signed(_T_885)}; // @[Parameters.scala 137:49]
  assign _T_888 = $signed(_T_886) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _T_889 = $signed(_T_888) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_890 = io_in_b_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31]
  assign _T_891 = {1'b0,$signed(_T_890)}; // @[Parameters.scala 137:49]
  assign _T_893 = $signed(_T_891) & -33'sh4000000; // @[Parameters.scala 137:52]
  assign _T_894 = $signed(_T_893) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_895 = io_in_b_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31]
  assign _T_896 = {1'b0,$signed(_T_895)}; // @[Parameters.scala 137:49]
  assign _T_898 = $signed(_T_896) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _T_899 = $signed(_T_898) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_903 = $signed(_T_868) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _T_904 = $signed(_T_903) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_905 = io_in_b_bits_address ^ 32'h10000; // @[Parameters.scala 137:31]
  assign _T_906 = {1'b0,$signed(_T_905)}; // @[Parameters.scala 137:49]
  assign _T_908 = $signed(_T_906) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _T_909 = $signed(_T_908) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_910 = io_in_b_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  assign _T_911 = {1'b0,$signed(_T_910)}; // @[Parameters.scala 137:49]
  assign _T_913 = $signed(_T_911) & -33'sh10000000; // @[Parameters.scala 137:52]
  assign _T_914 = $signed(_T_913) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_915 = io_in_b_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31]
  assign _T_916 = {1'b0,$signed(_T_915)}; // @[Parameters.scala 137:49]
  assign _T_918 = $signed(_T_916) & -33'sh20000000; // @[Parameters.scala 137:52]
  assign _T_919 = $signed(_T_918) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_921 = _T_889 | _T_894; // @[Parameters.scala 556:64]
  assign _T_922 = _T_921 | _T_899; // @[Parameters.scala 556:64]
  assign _T_923 = _T_922 | _T_904; // @[Parameters.scala 556:64]
  assign _T_924 = _T_923 | _T_909; // @[Parameters.scala 556:64]
  assign _T_925 = _T_924 | _T_914; // @[Parameters.scala 556:64]
  assign _T_926 = _T_925 | _T_919; // @[Parameters.scala 556:64]
  assign _T_928 = 27'hfff << io_in_b_bits_size; // @[package.scala 212:77]
  assign _GEN_72 = {{20'd0}, ~_T_928[11:0]}; // @[Edges.scala 22:16]
  assign _T_931 = io_in_b_bits_address & _GEN_72; // @[Edges.scala 22:16]
  assign _T_932 = _T_931 == 32'h0; // @[Edges.scala 22:24]
  assign _T_935 = 4'h1 << io_in_b_bits_size[1:0]; // @[OneHot.scala 65:12]
  assign _T_937 = _T_935[2:0] | 3'h1; // @[Misc.scala 201:81]
  assign _T_938 = io_in_b_bits_size >= 4'h3; // @[Misc.scala 205:21]
  assign _T_943 = _T_937[2] & ~io_in_b_bits_address[2]; // @[Misc.scala 214:38]
  assign _T_944 = _T_938 | _T_943; // @[Misc.scala 214:29]
  assign _T_946 = _T_937[2] & io_in_b_bits_address[2]; // @[Misc.scala 214:38]
  assign _T_947 = _T_938 | _T_946; // @[Misc.scala 214:29]
  assign _T_951 = ~io_in_b_bits_address[2] & ~io_in_b_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_952 = _T_937[1] & _T_951; // @[Misc.scala 214:38]
  assign _T_953 = _T_944 | _T_952; // @[Misc.scala 214:29]
  assign _T_954 = ~io_in_b_bits_address[2] & io_in_b_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_955 = _T_937[1] & _T_954; // @[Misc.scala 214:38]
  assign _T_956 = _T_944 | _T_955; // @[Misc.scala 214:29]
  assign _T_957 = io_in_b_bits_address[2] & ~io_in_b_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_958 = _T_937[1] & _T_957; // @[Misc.scala 214:38]
  assign _T_959 = _T_947 | _T_958; // @[Misc.scala 214:29]
  assign _T_960 = io_in_b_bits_address[2] & io_in_b_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_961 = _T_937[1] & _T_960; // @[Misc.scala 214:38]
  assign _T_962 = _T_947 | _T_961; // @[Misc.scala 214:29]
  assign _T_966 = _T_951 & ~io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_967 = _T_937[0] & _T_966; // @[Misc.scala 214:38]
  assign _T_968 = _T_953 | _T_967; // @[Misc.scala 214:29]
  assign _T_969 = _T_951 & io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_970 = _T_937[0] & _T_969; // @[Misc.scala 214:38]
  assign _T_971 = _T_953 | _T_970; // @[Misc.scala 214:29]
  assign _T_972 = _T_954 & ~io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_973 = _T_937[0] & _T_972; // @[Misc.scala 214:38]
  assign _T_974 = _T_956 | _T_973; // @[Misc.scala 214:29]
  assign _T_975 = _T_954 & io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_976 = _T_937[0] & _T_975; // @[Misc.scala 214:38]
  assign _T_977 = _T_956 | _T_976; // @[Misc.scala 214:29]
  assign _T_978 = _T_957 & ~io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_979 = _T_937[0] & _T_978; // @[Misc.scala 214:38]
  assign _T_980 = _T_959 | _T_979; // @[Misc.scala 214:29]
  assign _T_981 = _T_957 & io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_982 = _T_937[0] & _T_981; // @[Misc.scala 214:38]
  assign _T_983 = _T_959 | _T_982; // @[Misc.scala 214:29]
  assign _T_984 = _T_960 & ~io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_985 = _T_937[0] & _T_984; // @[Misc.scala 214:38]
  assign _T_986 = _T_962 | _T_985; // @[Misc.scala 214:29]
  assign _T_987 = _T_960 & io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_988 = _T_937[0] & _T_987; // @[Misc.scala 214:38]
  assign _T_989 = _T_962 | _T_988; // @[Misc.scala 214:29]
  assign _T_996 = {_T_989,_T_986,_T_983,_T_980,_T_977,_T_974,_T_971,_T_968}; // @[Cat.scala 29:58]
  assign _T_1004 = io_in_b_bits_source == io_in_b_bits_source; // @[Monitor.scala 165:113]
  assign _T_1005 = io_in_b_bits_opcode == 3'h6; // @[Monitor.scala 167:25]
  assign _T_1009 = 4'h6 == io_in_b_bits_size; // @[Parameters.scala 92:48]
  assign _T_1010 = ~io_in_b_bits_source & _T_1009; // @[Mux.scala 27:72]
  assign _T_1015 = io_in_b_bits_size <= 4'hc; // @[Parameters.scala 93:42]
  assign _T_1025 = _T_1010 & _T_1015; // @[Parameters.scala 1255:195]
  assign _T_1027 = _T_1025 | reset; // @[Monitor.scala 44:11]
  assign _T_1030 = _T_926 | reset; // @[Monitor.scala 44:11]
  assign _T_1033 = _T_1004 | reset; // @[Monitor.scala 44:11]
  assign _T_1036 = _T_932 | reset; // @[Monitor.scala 44:11]
  assign _T_1038 = io_in_b_bits_param <= 2'h2; // @[Bundles.scala 104:26]
  assign _T_1040 = _T_1038 | reset; // @[Monitor.scala 44:11]
  assign _T_1042 = io_in_b_bits_mask == _T_996; // @[Monitor.scala 173:30]
  assign _T_1044 = _T_1042 | reset; // @[Monitor.scala 44:11]
  assign _T_1048 = ~io_in_b_bits_corrupt | reset; // @[Monitor.scala 44:11]
  assign _T_1050 = io_in_b_bits_opcode == 3'h4; // @[Monitor.scala 177:25]
  assign _T_1075 = io_in_b_bits_param == 2'h0; // @[Monitor.scala 182:31]
  assign _T_1077 = _T_1075 | reset; // @[Monitor.scala 44:11]
  assign _T_1087 = io_in_b_bits_opcode == 3'h0; // @[Monitor.scala 187:25]
  assign _T_1120 = io_in_b_bits_opcode == 3'h1; // @[Monitor.scala 196:25]
  assign _T_1150 = io_in_b_bits_mask & ~_T_996; // @[Monitor.scala 202:31]
  assign _T_1151 = _T_1150 == 8'h0; // @[Monitor.scala 202:40]
  assign _T_1153 = _T_1151 | reset; // @[Monitor.scala 44:11]
  assign _T_1155 = io_in_b_bits_opcode == 3'h2; // @[Monitor.scala 205:25]
  assign _T_1188 = io_in_b_bits_opcode == 3'h3; // @[Monitor.scala 214:25]
  assign _T_1221 = io_in_b_bits_opcode == 3'h5; // @[Monitor.scala 223:25]
  assign _T_1261 = ~io_in_c_bits_source | io_in_c_bits_source; // @[Parameters.scala 1016:46]
  assign _T_1263 = 27'hfff << io_in_c_bits_size; // @[package.scala 212:77]
  assign _GEN_73 = {{20'd0}, ~_T_1263[11:0]}; // @[Edges.scala 22:16]
  assign _T_1266 = io_in_c_bits_address & _GEN_73; // @[Edges.scala 22:16]
  assign _T_1267 = _T_1266 == 32'h0; // @[Edges.scala 22:24]
  assign _T_1268 = io_in_c_bits_address ^ 32'h3000; // @[Parameters.scala 137:31]
  assign _T_1269 = {1'b0,$signed(_T_1268)}; // @[Parameters.scala 137:49]
  assign _T_1271 = $signed(_T_1269) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _T_1272 = $signed(_T_1271) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1273 = io_in_c_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31]
  assign _T_1274 = {1'b0,$signed(_T_1273)}; // @[Parameters.scala 137:49]
  assign _T_1276 = $signed(_T_1274) & -33'sh4000000; // @[Parameters.scala 137:52]
  assign _T_1277 = $signed(_T_1276) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1278 = io_in_c_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31]
  assign _T_1279 = {1'b0,$signed(_T_1278)}; // @[Parameters.scala 137:49]
  assign _T_1281 = $signed(_T_1279) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _T_1282 = $signed(_T_1281) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1284 = {1'b0,$signed(io_in_c_bits_address)}; // @[Parameters.scala 137:49]
  assign _T_1286 = $signed(_T_1284) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _T_1287 = $signed(_T_1286) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1288 = io_in_c_bits_address ^ 32'h10000; // @[Parameters.scala 137:31]
  assign _T_1289 = {1'b0,$signed(_T_1288)}; // @[Parameters.scala 137:49]
  assign _T_1291 = $signed(_T_1289) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _T_1292 = $signed(_T_1291) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1293 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  assign _T_1294 = {1'b0,$signed(_T_1293)}; // @[Parameters.scala 137:49]
  assign _T_1296 = $signed(_T_1294) & -33'sh10000000; // @[Parameters.scala 137:52]
  assign _T_1297 = $signed(_T_1296) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1298 = io_in_c_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31]
  assign _T_1299 = {1'b0,$signed(_T_1298)}; // @[Parameters.scala 137:49]
  assign _T_1301 = $signed(_T_1299) & -33'sh20000000; // @[Parameters.scala 137:52]
  assign _T_1302 = $signed(_T_1301) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1304 = _T_1272 | _T_1277; // @[Parameters.scala 556:64]
  assign _T_1305 = _T_1304 | _T_1282; // @[Parameters.scala 556:64]
  assign _T_1306 = _T_1305 | _T_1287; // @[Parameters.scala 556:64]
  assign _T_1307 = _T_1306 | _T_1292; // @[Parameters.scala 556:64]
  assign _T_1308 = _T_1307 | _T_1297; // @[Parameters.scala 556:64]
  assign _T_1309 = _T_1308 | _T_1302; // @[Parameters.scala 556:64]
  assign _T_1330 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 242:25]
  assign _T_1332 = _T_1309 | reset; // @[Monitor.scala 44:11]
  assign _T_1335 = _T_1261 | reset; // @[Monitor.scala 44:11]
  assign _T_1337 = io_in_c_bits_size >= 4'h3; // @[Monitor.scala 245:30]
  assign _T_1339 = _T_1337 | reset; // @[Monitor.scala 44:11]
  assign _T_1342 = _T_1267 | reset; // @[Monitor.scala 44:11]
  assign _T_1344 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 122:29]
  assign _T_1346 = _T_1344 | reset; // @[Monitor.scala 44:11]
  assign _T_1352 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 251:25]
  assign _T_1370 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 259:25]
  assign _T_1372 = io_in_c_bits_size <= 4'hc; // @[Parameters.scala 93:42]
  assign _T_1377 = _T_1372 & _T_1261; // @[Parameters.scala 1066:30]
  assign _T_1387 = io_in_c_bits_size <= 4'h6; // @[Parameters.scala 93:42]
  assign _T_1393 = $signed(_T_1294) & 33'sh80000000; // @[Parameters.scala 137:52]
  assign _T_1394 = $signed(_T_1393) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1395 = _T_1387 & _T_1394; // @[Parameters.scala 601:56]
  assign _T_1398 = _T_1377 & _T_1395; // @[Parameters.scala 1240:195]
  assign _T_1400 = _T_1398 | reset; // @[Monitor.scala 44:11]
  assign _T_1405 = 4'h6 == io_in_c_bits_size; // @[Parameters.scala 92:48]
  assign _T_1406 = ~io_in_c_bits_source & _T_1405; // @[Mux.scala 27:72]
  assign _T_1421 = _T_1406 & _T_1372; // @[Parameters.scala 1255:195]
  assign _T_1423 = _T_1421 | reset; // @[Monitor.scala 44:11]
  assign _T_1435 = io_in_c_bits_param <= 3'h2; // @[Bundles.scala 116:29]
  assign _T_1437 = _T_1435 | reset; // @[Monitor.scala 44:11]
  assign _T_1443 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 269:25]
  assign _T_1512 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 278:25]
  assign _T_1522 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 282:31]
  assign _T_1524 = _T_1522 | reset; // @[Monitor.scala 44:11]
  assign _T_1530 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 286:25]
  assign _T_1544 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 293:25]
  assign _T_1566 = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  assign _T_1571 = ~_T_9[11:3]; // @[Edges.scala 221:59]
  assign _T_1577 = _T_1575 - 9'h1; // @[Edges.scala 231:28]
  assign _T_1578 = _T_1575 == 9'h0; // @[Edges.scala 232:25]
  assign _T_1592 = io_in_a_valid & ~_T_1578; // @[Monitor.scala 389:19]
  assign _T_1593 = io_in_a_bits_opcode == _T_1586; // @[Monitor.scala 390:32]
  assign _T_1595 = _T_1593 | reset; // @[Monitor.scala 44:11]
  assign _T_1597 = io_in_a_bits_param == _T_1587; // @[Monitor.scala 391:32]
  assign _T_1599 = _T_1597 | reset; // @[Monitor.scala 44:11]
  assign _T_1601 = io_in_a_bits_size == _T_1588; // @[Monitor.scala 392:32]
  assign _T_1603 = _T_1601 | reset; // @[Monitor.scala 44:11]
  assign _T_1605 = io_in_a_bits_source == _T_1589; // @[Monitor.scala 393:32]
  assign _T_1607 = _T_1605 | reset; // @[Monitor.scala 44:11]
  assign _T_1609 = io_in_a_bits_address == _T_1590; // @[Monitor.scala 394:32]
  assign _T_1611 = _T_1609 | reset; // @[Monitor.scala 44:11]
  assign _T_1614 = _T_1566 & _T_1578; // @[Monitor.scala 396:20]
  assign _T_1615 = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  assign _T_1617 = 27'hfff << io_in_d_bits_size; // @[package.scala 212:77]
  assign _T_1620 = ~_T_1617[11:3]; // @[Edges.scala 221:59]
  assign _T_1625 = _T_1623 - 9'h1; // @[Edges.scala 231:28]
  assign _T_1626 = _T_1623 == 9'h0; // @[Edges.scala 232:25]
  assign _T_1641 = io_in_d_valid & ~_T_1626; // @[Monitor.scala 541:19]
  assign _T_1642 = io_in_d_bits_opcode == _T_1634; // @[Monitor.scala 542:29]
  assign _T_1644 = _T_1642 | reset; // @[Monitor.scala 51:11]
  assign _T_1646 = io_in_d_bits_param == _T_1635; // @[Monitor.scala 543:29]
  assign _T_1648 = _T_1646 | reset; // @[Monitor.scala 51:11]
  assign _T_1650 = io_in_d_bits_size == _T_1636; // @[Monitor.scala 544:29]
  assign _T_1652 = _T_1650 | reset; // @[Monitor.scala 51:11]
  assign _T_1654 = io_in_d_bits_source == _T_1637; // @[Monitor.scala 545:29]
  assign _T_1656 = _T_1654 | reset; // @[Monitor.scala 51:11]
  assign _T_1658 = io_in_d_bits_sink == _T_1638; // @[Monitor.scala 546:29]
  assign _T_1660 = _T_1658 | reset; // @[Monitor.scala 51:11]
  assign _T_1662 = io_in_d_bits_denied == _T_1639; // @[Monitor.scala 547:29]
  assign _T_1664 = _T_1662 | reset; // @[Monitor.scala 51:11]
  assign _T_1667 = _T_1615 & _T_1626; // @[Monitor.scala 549:20]
  assign _T_1668 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37]
  assign _T_1679 = _T_1677 - 9'h1; // @[Edges.scala 231:28]
  assign _T_1680 = _T_1677 == 9'h0; // @[Edges.scala 232:25]
  assign _T_1694 = io_in_b_valid & ~_T_1680; // @[Monitor.scala 412:19]
  assign _T_1695 = io_in_b_bits_opcode == _T_1688; // @[Monitor.scala 413:32]
  assign _T_1697 = _T_1695 | reset; // @[Monitor.scala 44:11]
  assign _T_1699 = io_in_b_bits_param == _T_1689; // @[Monitor.scala 414:32]
  assign _T_1701 = _T_1699 | reset; // @[Monitor.scala 44:11]
  assign _T_1703 = io_in_b_bits_size == _T_1690; // @[Monitor.scala 415:32]
  assign _T_1705 = _T_1703 | reset; // @[Monitor.scala 44:11]
  assign _T_1707 = io_in_b_bits_source == _T_1691; // @[Monitor.scala 416:32]
  assign _T_1709 = _T_1707 | reset; // @[Monitor.scala 44:11]
  assign _T_1711 = io_in_b_bits_address == _T_1692; // @[Monitor.scala 417:32]
  assign _T_1713 = _T_1711 | reset; // @[Monitor.scala 44:11]
  assign _T_1716 = _T_1668 & _T_1680; // @[Monitor.scala 419:20]
  assign _T_1717 = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37]
  assign _T_1722 = ~_T_1263[11:3]; // @[Edges.scala 221:59]
  assign _T_1727 = _T_1725 - 9'h1; // @[Edges.scala 231:28]
  assign _T_1728 = _T_1725 == 9'h0; // @[Edges.scala 232:25]
  assign _T_1742 = io_in_c_valid & ~_T_1728; // @[Monitor.scala 517:19]
  assign _T_1743 = io_in_c_bits_opcode == _T_1736; // @[Monitor.scala 518:32]
  assign _T_1745 = _T_1743 | reset; // @[Monitor.scala 44:11]
  assign _T_1747 = io_in_c_bits_param == _T_1737; // @[Monitor.scala 519:32]
  assign _T_1749 = _T_1747 | reset; // @[Monitor.scala 44:11]
  assign _T_1751 = io_in_c_bits_size == _T_1738; // @[Monitor.scala 520:32]
  assign _T_1753 = _T_1751 | reset; // @[Monitor.scala 44:11]
  assign _T_1755 = io_in_c_bits_source == _T_1739; // @[Monitor.scala 521:32]
  assign _T_1757 = _T_1755 | reset; // @[Monitor.scala 44:11]
  assign _T_1759 = io_in_c_bits_address == _T_1740; // @[Monitor.scala 522:32]
  assign _T_1761 = _T_1759 | reset; // @[Monitor.scala 44:11]
  assign _T_1764 = _T_1717 & _T_1728; // @[Monitor.scala 524:20]
  assign _T_1776 = _T_1774 - 9'h1; // @[Edges.scala 231:28]
  assign a_first = _T_1774 == 9'h0; // @[Edges.scala 232:25]
  assign _T_1794 = _T_1792 - 9'h1; // @[Edges.scala 231:28]
  assign d_first = _T_1792 == 9'h0; // @[Edges.scala 232:25]
  assign _GEN_74 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 632:69]
  assign _T_1802 = {{1'd0}, _GEN_74}; // @[Monitor.scala 632:69]
  assign _T_1803 = inflight_opcodes >> _T_1802; // @[Monitor.scala 632:44]
  assign _T_1807 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  assign _GEN_75 = {{8'd0}, _T_1803}; // @[Monitor.scala 632:97]
  assign _T_1808 = _GEN_75 & _T_1807; // @[Monitor.scala 632:97]
  assign _T_1809 = {{1'd0}, _T_1808[15:1]}; // @[Monitor.scala 632:152]
  assign _T_1810 = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 636:65]
  assign _T_1811 = inflight_sizes >> _T_1810; // @[Monitor.scala 636:40]
  assign _T_1815 = 16'h100 - 16'h1; // @[Monitor.scala 609:57]
  assign _T_1816 = _T_1811 & _T_1815; // @[Monitor.scala 636:91]
  assign _T_1817 = {{1'd0}, _T_1816[15:1]}; // @[Monitor.scala 636:144]
  assign _T_1821 = _T_1566 & a_first; // @[Monitor.scala 646:27]
  assign _T_1823 = 2'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  assign _T_1824 = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 648:53]
  assign _T_1825 = _T_1824 | 4'h1; // @[Monitor.scala 648:61]
  assign _T_1826 = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 649:49]
  assign _T_1827 = _T_1826 | 5'h1; // @[Monitor.scala 649:57]
  assign _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 650:72]
  assign _T_1828 = {{1'd0}, _GEN_78}; // @[Monitor.scala 650:72]
  assign a_opcodes_set_interm = _T_1821 ? _T_1825 : 4'h0; // @[Monitor.scala 646:72]
  assign _GEN_79 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 650:47]
  assign _T_1829 = _GEN_79 << _T_1828; // @[Monitor.scala 650:47]
  assign _T_1830 = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 651:68]
  assign a_sizes_set_interm = _T_1821 ? _T_1827 : 5'h0; // @[Monitor.scala 646:72]
  assign _GEN_80 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 651:43]
  assign _T_1831 = _GEN_80 << _T_1830; // @[Monitor.scala 651:43]
  assign _T_1832 = inflight >> io_in_a_bits_source; // @[Monitor.scala 652:26]
  assign _T_1836 = ~_T_1832[0] | reset; // @[Monitor.scala 44:11]
  assign a_set = _T_1821 ? _T_1823 : 2'h0; // @[Monitor.scala 646:72]
  assign _GEN_30 = _T_1821 ? _T_1829 : 19'h0; // @[Monitor.scala 646:72]
  assign _GEN_31 = _T_1821 ? _T_1831 : 20'h0; // @[Monitor.scala 646:72]
  assign _T_1840 = _T_1615 & d_first; // @[Monitor.scala 663:27]
  assign _T_1843 = _T_1840 & ~_T_732; // @[Monitor.scala 663:72]
  assign _T_1844 = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  assign _GEN_82 = {{15'd0}, _T_1807}; // @[Monitor.scala 665:76]
  assign _T_1850 = _GEN_82 << _T_1802; // @[Monitor.scala 665:76]
  assign _GEN_83 = {{15'd0}, _T_1815}; // @[Monitor.scala 666:72]
  assign _T_1856 = _GEN_83 << _T_1810; // @[Monitor.scala 666:72]
  assign d_clr = _T_1843 ? _T_1844 : 2'h0; // @[Monitor.scala 663:91]
  assign _GEN_33 = _T_1843 ? _T_1850 : 31'h0; // @[Monitor.scala 663:91]
  assign _GEN_34 = _T_1843 ? _T_1856 : 31'h0; // @[Monitor.scala 663:91]
  assign _T_1857 = io_in_d_valid & d_first; // @[Monitor.scala 668:26]
  assign _T_1860 = _T_1857 & ~_T_732; // @[Monitor.scala 668:71]
  assign _T_1861 = inflight >> io_in_d_bits_source; // @[Monitor.scala 669:25]
  assign _T_1863 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 669:93]
  assign _T_1864 = io_in_a_valid & _T_1863; // @[Monitor.scala 669:68]
  assign _T_1865 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 669:142]
  assign _T_1866 = _T_1864 & _T_1865; // @[Monitor.scala 669:119]
  assign _T_1867 = _T_1866 & a_first; // @[Monitor.scala 669:166]
  assign _T_1868 = _T_1861[0] | _T_1867; // @[Monitor.scala 669:49]
  assign _T_1870 = _T_1868 | reset; // @[Monitor.scala 51:11]
  assign a_opcode_lookup = _T_1809[3:0]; // @[Monitor.scala 632:21]
  assign _GEN_37 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 670:37]
  assign _GEN_38 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_37; // @[Monitor.scala 670:37]
  assign _GEN_39 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_38; // @[Monitor.scala 670:37]
  assign _GEN_40 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_39; // @[Monitor.scala 670:37]
  assign _GEN_41 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_40; // @[Monitor.scala 670:37]
  assign _GEN_42 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_41; // @[Monitor.scala 670:37]
  assign _T_1873 = io_in_d_bits_opcode == _GEN_42; // @[Monitor.scala 670:37]
  assign _GEN_49 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_40; // @[Monitor.scala 670:96]
  assign _GEN_50 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_49; // @[Monitor.scala 670:96]
  assign _T_1875 = io_in_d_bits_opcode == _GEN_50; // @[Monitor.scala 670:96]
  assign _T_1876 = _T_1873 | _T_1875; // @[Monitor.scala 670:71]
  assign _GEN_53 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 671:60]
  assign _GEN_54 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_53; // @[Monitor.scala 671:60]
  assign _GEN_55 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_54; // @[Monitor.scala 671:60]
  assign _GEN_56 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_55; // @[Monitor.scala 671:60]
  assign _GEN_57 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_56; // @[Monitor.scala 671:60]
  assign _GEN_58 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_57; // @[Monitor.scala 671:60]
  assign _T_1877 = io_in_d_bits_opcode == _GEN_58; // @[Monitor.scala 671:60]
  assign _GEN_65 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_56; // @[Monitor.scala 671:124]
  assign _GEN_66 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_65; // @[Monitor.scala 671:124]
  assign _T_1878 = io_in_d_bits_opcode == _GEN_66; // @[Monitor.scala 671:124]
  assign _T_1879 = _T_1877 | _T_1878; // @[Monitor.scala 671:99]
  assign _T_1880 = io_in_a_valid & _T_1879; // @[Monitor.scala 671:34]
  assign _T_1881 = _T_1876 | _T_1880; // @[Monitor.scala 671:15]
  assign _T_1883 = _T_1881 | reset; // @[Monitor.scala 51:11]
  assign a_size_lookup = _T_1817[7:0]; // @[Monitor.scala 636:19]
  assign _GEN_84 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 673:34]
  assign _T_1885 = _GEN_84 == a_size_lookup; // @[Monitor.scala 673:34]
  assign _T_1887 = io_in_a_valid & _T_1865; // @[Monitor.scala 673:72]
  assign _T_1888 = _T_1885 | _T_1887; // @[Monitor.scala 673:53]
  assign _T_1890 = _T_1888 | reset; // @[Monitor.scala 51:11]
  assign _T_1893 = _T_1857 & a_first; // @[Monitor.scala 675:36]
  assign _T_1894 = _T_1893 & io_in_a_valid; // @[Monitor.scala 675:47]
  assign _T_1896 = _T_1894 & _T_1863; // @[Monitor.scala 675:65]
  assign _T_1898 = _T_1896 & ~_T_732; // @[Monitor.scala 675:116]
  assign _T_1900 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 676:32]
  assign _T_1902 = _T_1900 | reset; // @[Monitor.scala 51:11]
  assign _T_1904 = a_set != d_clr; // @[Monitor.scala 680:20]
  assign _T_1905 = |a_set; // @[Monitor.scala 680:40]
  assign _T_1907 = _T_1904 | ~_T_1905; // @[Monitor.scala 680:30]
  assign _T_1909 = _T_1907 | reset; // @[Monitor.scala 51:11]
  assign _T_1911 = inflight | a_set; // @[Monitor.scala 683:27]
  assign _T_1913 = _T_1911 & ~d_clr; // @[Monitor.scala 683:36]
  assign a_opcodes_set = _GEN_30[7:0]; // @[Monitor.scala 650:21]
  assign _T_1914 = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 684:43]
  assign d_opcodes_clr = _GEN_33[7:0]; // @[Monitor.scala 665:21]
  assign _T_1916 = _T_1914 & ~d_opcodes_clr; // @[Monitor.scala 684:60]
  assign a_sizes_set = _GEN_31[15:0]; // @[Monitor.scala 651:19]
  assign _T_1917 = inflight_sizes | a_sizes_set; // @[Monitor.scala 685:39]
  assign d_sizes_clr = _GEN_34[15:0]; // @[Monitor.scala 666:19]
  assign _T_1919 = _T_1917 & ~d_sizes_clr; // @[Monitor.scala 685:54]
  assign _T_1946 = _T_1944 - 9'h1; // @[Edges.scala 231:28]
  assign _T_1947 = _T_1944 == 9'h0; // @[Edges.scala 232:25]
  assign _T_1957 = _T_1615 & _T_1947; // @[Monitor.scala 703:27]
  assign _T_1961 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 72:40]
  assign _T_1962 = _T_1957 & _T_1961; // @[Monitor.scala 703:38]
  assign _T_1963 = 4'h1 << io_in_d_bits_sink; // @[OneHot.scala 58:35]
  assign _T_1964 = _T_1935 >> io_in_d_bits_sink; // @[Monitor.scala 705:23]
  assign _T_1968 = ~_T_1964[0] | reset; // @[Monitor.scala 51:11]
  assign _GEN_69 = _T_1962 ? _T_1963 : 4'h0; // @[Monitor.scala 703:72]
  assign _T_1971 = io_in_e_ready & io_in_e_valid; // @[Decoupled.scala 40:37]
  assign _T_1974 = 4'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35]
  assign _T_1975 = _GEN_69 | _T_1935; // @[Monitor.scala 711:24]
  assign _T_1976 = _T_1975 >> io_in_e_bits_sink; // @[Monitor.scala 711:35]
  assign _T_1979 = _T_1976[0] | reset; // @[Monitor.scala 44:11]
  assign _GEN_70 = _T_1971 ? _T_1974 : 4'h0; // @[Monitor.scala 709:73]
  assign _T_1981 = _T_1935 | _GEN_69; // @[Monitor.scala 716:27]
  assign _T_1983 = _T_1981 & ~_GEN_70; // @[Monitor.scala 716:36]
  assign _GEN_85 = io_in_a_valid & _T_98; // @[Monitor.scala 44:11]
  assign _GEN_99 = io_in_a_valid & _T_176; // @[Monitor.scala 44:11]
  assign _GEN_115 = io_in_a_valid & _T_258; // @[Monitor.scala 44:11]
  assign _GEN_125 = io_in_a_valid & _T_341; // @[Monitor.scala 44:11]
  assign _GEN_135 = io_in_a_valid & _T_427; // @[Monitor.scala 44:11]
  assign _GEN_145 = io_in_a_valid & _T_515; // @[Monitor.scala 44:11]
  assign _GEN_155 = io_in_a_valid & _T_579; // @[Monitor.scala 44:11]
  assign _GEN_165 = io_in_a_valid & _T_643; // @[Monitor.scala 44:11]
  assign _GEN_175 = io_in_d_valid & _T_732; // @[Monitor.scala 51:11]
  assign _GEN_185 = io_in_d_valid & _T_752; // @[Monitor.scala 51:11]
  assign _GEN_195 = io_in_d_valid & _T_780; // @[Monitor.scala 51:11]
  assign _GEN_205 = io_in_d_valid & _T_809; // @[Monitor.scala 51:11]
  assign _GEN_211 = io_in_d_valid & _T_826; // @[Monitor.scala 51:11]
  assign _GEN_217 = io_in_d_valid & _T_844; // @[Monitor.scala 51:11]
  assign _GEN_223 = io_in_b_valid & _T_1005; // @[Monitor.scala 44:11]
  assign _GEN_237 = io_in_b_valid & _T_1050; // @[Monitor.scala 44:11]
  assign _GEN_251 = io_in_b_valid & _T_1087; // @[Monitor.scala 44:11]
  assign _GEN_263 = io_in_b_valid & _T_1120; // @[Monitor.scala 44:11]
  assign _GEN_275 = io_in_b_valid & _T_1155; // @[Monitor.scala 44:11]
  assign _GEN_285 = io_in_b_valid & _T_1188; // @[Monitor.scala 44:11]
  assign _GEN_295 = io_in_b_valid & _T_1221; // @[Monitor.scala 44:11]
  assign _GEN_307 = io_in_c_valid & _T_1330; // @[Monitor.scala 44:11]
  assign _GEN_317 = io_in_c_valid & _T_1352; // @[Monitor.scala 44:11]
  assign _GEN_327 = io_in_c_valid & _T_1370; // @[Monitor.scala 44:11]
  assign _GEN_339 = io_in_c_valid & _T_1443; // @[Monitor.scala 44:11]
  assign _GEN_351 = io_in_c_valid & _T_1512; // @[Monitor.scala 44:11]
  assign _GEN_359 = io_in_c_valid & _T_1530; // @[Monitor.scala 44:11]
  assign _GEN_367 = io_in_c_valid & _T_1544; // @[Monitor.scala 44:11]
  assign TLMonitor_35_covSum = 30'h0;
  assign io_covSum = TLMonitor_35_covSum;
  assign stopEn0 = _GEN_85 & ~_T_128;
  assign stopEn1 = _GEN_85 & ~_T_151;
  assign stopEn2 = _GEN_85 & ~_T_154;
  assign stopEn3 = _GEN_85 & ~_T_158;
  assign stopEn4 = _GEN_85 & ~_T_161;
  assign stopEn5 = _GEN_85 & ~_T_165;
  assign stopEn6 = _GEN_85 & ~_T_170;
  assign stopEn7 = _GEN_99 & ~_T_128;
  assign stopEn8 = _GEN_99 & ~_T_151;
  assign stopEn9 = _GEN_99 & ~_T_154;
  assign stopEn10 = _GEN_99 & ~_T_158;
  assign stopEn11 = _GEN_99 & ~_T_161;
  assign stopEn12 = _GEN_99 & ~_T_165;
  assign stopEn13 = _GEN_99 & ~_T_247;
  assign stopEn14 = _GEN_99 & ~_T_170;
  assign stopEn15 = _GEN_115 & ~_T_321;
  assign stopEn16 = _GEN_115 & ~_T_154;
  assign stopEn17 = _GEN_115 & ~_T_161;
  assign stopEn18 = _GEN_115 & ~_T_331;
  assign stopEn19 = _GEN_115 & ~_T_335;
  assign stopEn20 = _GEN_125 & ~_T_411;
  assign stopEn21 = _GEN_125 & ~_T_154;
  assign stopEn22 = _GEN_125 & ~_T_161;
  assign stopEn23 = _GEN_125 & ~_T_331;
  assign stopEn24 = _GEN_125 & ~_T_335;
  assign stopEn25 = _GEN_135 & ~_T_411;
  assign stopEn26 = _GEN_135 & ~_T_154;
  assign stopEn27 = _GEN_135 & ~_T_161;
  assign stopEn28 = _GEN_135 & ~_T_331;
  assign stopEn29 = _GEN_135 & ~_T_513;
  assign stopEn30 = _GEN_145 & ~_T_563;
  assign stopEn31 = _GEN_145 & ~_T_154;
  assign stopEn32 = _GEN_145 & ~_T_161;
  assign stopEn33 = _GEN_145 & ~_T_573;
  assign stopEn34 = _GEN_145 & ~_T_335;
  assign stopEn35 = _GEN_155 & ~_T_563;
  assign stopEn36 = _GEN_155 & ~_T_154;
  assign stopEn37 = _GEN_155 & ~_T_161;
  assign stopEn38 = _GEN_155 & ~_T_637;
  assign stopEn39 = _GEN_155 & ~_T_335;
  assign stopEn40 = _GEN_165 & ~_T_703;
  assign stopEn41 = _GEN_165 & ~_T_154;
  assign stopEn42 = _GEN_165 & ~_T_161;
  assign stopEn43 = _GEN_165 & ~_T_713;
  assign stopEn44 = _GEN_165 & ~_T_335;
  assign stopEn45 = io_in_d_valid & ~_T_725;
  assign stopEn46 = _GEN_175 & ~_T_734;
  assign stopEn47 = _GEN_175 & ~_T_738;
  assign stopEn48 = _GEN_175 & ~_T_742;
  assign stopEn49 = _GEN_175 & ~_T_746;
  assign stopEn50 = _GEN_175 & ~_T_750;
  assign stopEn51 = _GEN_185 & ~_T_734;
  assign stopEn52 = _GEN_185 & ~_T_738;
  assign stopEn53 = _GEN_185 & ~_T_765;
  assign stopEn54 = _GEN_185 & ~_T_769;
  assign stopEn55 = _GEN_185 & ~_T_746;
  assign stopEn56 = _GEN_195 & ~_T_734;
  assign stopEn57 = _GEN_195 & ~_T_738;
  assign stopEn58 = _GEN_195 & ~_T_765;
  assign stopEn59 = _GEN_195 & ~_T_769;
  assign stopEn60 = _GEN_195 & ~_T_802;
  assign stopEn61 = _GEN_205 & ~_T_734;
  assign stopEn62 = _GEN_205 & ~_T_742;
  assign stopEn63 = _GEN_205 & ~_T_746;
  assign stopEn64 = _GEN_211 & ~_T_734;
  assign stopEn65 = _GEN_211 & ~_T_742;
  assign stopEn66 = _GEN_211 & ~_T_802;
  assign stopEn67 = _GEN_217 & ~_T_734;
  assign stopEn68 = _GEN_217 & ~_T_742;
  assign stopEn69 = _GEN_217 & ~_T_746;
  assign stopEn70 = io_in_b_valid & ~_T_863;
  assign stopEn71 = _GEN_223 & ~_T_1027;
  assign stopEn72 = _GEN_223 & ~_T_1030;
  assign stopEn73 = _GEN_223 & ~_T_1033;
  assign stopEn74 = _GEN_223 & ~_T_1036;
  assign stopEn75 = _GEN_223 & ~_T_1040;
  assign stopEn76 = _GEN_223 & ~_T_1044;
  assign stopEn77 = _GEN_223 & ~_T_1048;
  assign stopEn78 = _GEN_237 & ~reset;
  assign stopEn79 = _GEN_237 & ~_T_1030;
  assign stopEn80 = _GEN_237 & ~_T_1033;
  assign stopEn81 = _GEN_237 & ~_T_1036;
  assign stopEn82 = _GEN_237 & ~_T_1077;
  assign stopEn83 = _GEN_237 & ~_T_1044;
  assign stopEn84 = _GEN_237 & ~_T_1048;
  assign stopEn85 = _GEN_251 & ~reset;
  assign stopEn86 = _GEN_251 & ~_T_1030;
  assign stopEn87 = _GEN_251 & ~_T_1033;
  assign stopEn88 = _GEN_251 & ~_T_1036;
  assign stopEn89 = _GEN_251 & ~_T_1077;
  assign stopEn90 = _GEN_251 & ~_T_1044;
  assign stopEn91 = _GEN_263 & ~reset;
  assign stopEn92 = _GEN_263 & ~_T_1030;
  assign stopEn93 = _GEN_263 & ~_T_1033;
  assign stopEn94 = _GEN_263 & ~_T_1036;
  assign stopEn95 = _GEN_263 & ~_T_1077;
  assign stopEn96 = _GEN_263 & ~_T_1153;
  assign stopEn97 = _GEN_275 & ~reset;
  assign stopEn98 = _GEN_275 & ~_T_1030;
  assign stopEn99 = _GEN_275 & ~_T_1033;
  assign stopEn100 = _GEN_275 & ~_T_1036;
  assign stopEn101 = _GEN_275 & ~_T_1044;
  assign stopEn102 = _GEN_285 & ~reset;
  assign stopEn103 = _GEN_285 & ~_T_1030;
  assign stopEn104 = _GEN_285 & ~_T_1033;
  assign stopEn105 = _GEN_285 & ~_T_1036;
  assign stopEn106 = _GEN_285 & ~_T_1044;
  assign stopEn107 = _GEN_295 & ~reset;
  assign stopEn108 = _GEN_295 & ~_T_1030;
  assign stopEn109 = _GEN_295 & ~_T_1033;
  assign stopEn110 = _GEN_295 & ~_T_1036;
  assign stopEn111 = _GEN_295 & ~_T_1044;
  assign stopEn112 = _GEN_295 & ~_T_1048;
  assign stopEn113 = _GEN_307 & ~_T_1332;
  assign stopEn114 = _GEN_307 & ~_T_1335;
  assign stopEn115 = _GEN_307 & ~_T_1339;
  assign stopEn116 = _GEN_307 & ~_T_1342;
  assign stopEn117 = _GEN_307 & ~_T_1346;
  assign stopEn118 = _GEN_317 & ~_T_1332;
  assign stopEn119 = _GEN_317 & ~_T_1335;
  assign stopEn120 = _GEN_317 & ~_T_1339;
  assign stopEn121 = _GEN_317 & ~_T_1342;
  assign stopEn122 = _GEN_317 & ~_T_1346;
  assign stopEn123 = _GEN_327 & ~_T_1400;
  assign stopEn124 = _GEN_327 & ~_T_1423;
  assign stopEn125 = _GEN_327 & ~_T_1335;
  assign stopEn126 = _GEN_327 & ~_T_1339;
  assign stopEn127 = _GEN_327 & ~_T_1342;
  assign stopEn128 = _GEN_327 & ~_T_1437;
  assign stopEn129 = _GEN_339 & ~_T_1400;
  assign stopEn130 = _GEN_339 & ~_T_1423;
  assign stopEn131 = _GEN_339 & ~_T_1335;
  assign stopEn132 = _GEN_339 & ~_T_1339;
  assign stopEn133 = _GEN_339 & ~_T_1342;
  assign stopEn134 = _GEN_339 & ~_T_1437;
  assign stopEn135 = _GEN_351 & ~_T_1332;
  assign stopEn136 = _GEN_351 & ~_T_1335;
  assign stopEn137 = _GEN_351 & ~_T_1342;
  assign stopEn138 = _GEN_351 & ~_T_1524;
  assign stopEn139 = _GEN_359 & ~_T_1332;
  assign stopEn140 = _GEN_359 & ~_T_1335;
  assign stopEn141 = _GEN_359 & ~_T_1342;
  assign stopEn142 = _GEN_359 & ~_T_1524;
  assign stopEn143 = _GEN_367 & ~_T_1332;
  assign stopEn144 = _GEN_367 & ~_T_1335;
  assign stopEn145 = _GEN_367 & ~_T_1342;
  assign stopEn146 = _GEN_367 & ~_T_1524;
  assign stopEn147 = _T_1592 & ~_T_1595;
  assign stopEn148 = _T_1592 & ~_T_1599;
  assign stopEn149 = _T_1592 & ~_T_1603;
  assign stopEn150 = _T_1592 & ~_T_1607;
  assign stopEn151 = _T_1592 & ~_T_1611;
  assign stopEn152 = _T_1641 & ~_T_1644;
  assign stopEn153 = _T_1641 & ~_T_1648;
  assign stopEn154 = _T_1641 & ~_T_1652;
  assign stopEn155 = _T_1641 & ~_T_1656;
  assign stopEn156 = _T_1641 & ~_T_1660;
  assign stopEn157 = _T_1641 & ~_T_1664;
  assign stopEn158 = _T_1694 & ~_T_1697;
  assign stopEn159 = _T_1694 & ~_T_1701;
  assign stopEn160 = _T_1694 & ~_T_1705;
  assign stopEn161 = _T_1694 & ~_T_1709;
  assign stopEn162 = _T_1694 & ~_T_1713;
  assign stopEn163 = _T_1742 & ~_T_1745;
  assign stopEn164 = _T_1742 & ~_T_1749;
  assign stopEn165 = _T_1742 & ~_T_1753;
  assign stopEn166 = _T_1742 & ~_T_1757;
  assign stopEn167 = _T_1742 & ~_T_1761;
  assign stopEn168 = _T_1821 & ~_T_1836;
  assign stopEn169 = _T_1860 & ~_T_1870;
  assign stopEn170 = _T_1860 & ~_T_1883;
  assign stopEn171 = _T_1860 & ~_T_1890;
  assign stopEn172 = _T_1898 & ~_T_1902;
  assign stopEn173 = ~_T_1909;
  assign stopEn174 = _T_1962 & ~_T_1968;
  assign stopEn175 = _T_1971 & ~_T_1979;
  assign TLMonitor_35_or63 = stopEn0 | stopEn1;
  assign TLMonitor_35_or130 = stopEn3 | stopEn4;
  assign TLMonitor_35_or64 = stopEn2 | TLMonitor_35_or130;
  assign TLMonitor_35_or31 = TLMonitor_35_or63 | TLMonitor_35_or64;
  assign TLMonitor_35_or132 = stopEn6 | stopEn7;
  assign TLMonitor_35_or65 = stopEn5 | TLMonitor_35_or132;
  assign TLMonitor_35_or134 = stopEn9 | stopEn10;
  assign TLMonitor_35_or66 = stopEn8 | TLMonitor_35_or134;
  assign TLMonitor_35_or32 = TLMonitor_35_or65 | TLMonitor_35_or66;
  assign TLMonitor_35_or15 = TLMonitor_35_or31 | TLMonitor_35_or32;
  assign TLMonitor_35_or67 = stopEn11 | stopEn12;
  assign TLMonitor_35_or138 = stopEn14 | stopEn15;
  assign TLMonitor_35_or68 = stopEn13 | TLMonitor_35_or138;
  assign TLMonitor_35_or33 = TLMonitor_35_or67 | TLMonitor_35_or68;
  assign TLMonitor_35_or140 = stopEn17 | stopEn18;
  assign TLMonitor_35_or69 = stopEn16 | TLMonitor_35_or140;
  assign TLMonitor_35_or142 = stopEn20 | stopEn21;
  assign TLMonitor_35_or70 = stopEn19 | TLMonitor_35_or142;
  assign TLMonitor_35_or34 = TLMonitor_35_or69 | TLMonitor_35_or70;
  assign TLMonitor_35_or16 = TLMonitor_35_or33 | TLMonitor_35_or34;
  assign TLMonitor_35_or7 = TLMonitor_35_or15 | TLMonitor_35_or16;
  assign TLMonitor_35_or71 = stopEn22 | stopEn23;
  assign TLMonitor_35_or146 = stopEn25 | stopEn26;
  assign TLMonitor_35_or72 = stopEn24 | TLMonitor_35_or146;
  assign TLMonitor_35_or35 = TLMonitor_35_or71 | TLMonitor_35_or72;
  assign TLMonitor_35_or148 = stopEn28 | stopEn29;
  assign TLMonitor_35_or73 = stopEn27 | TLMonitor_35_or148;
  assign TLMonitor_35_or150 = stopEn31 | stopEn32;
  assign TLMonitor_35_or74 = stopEn30 | TLMonitor_35_or150;
  assign TLMonitor_35_or36 = TLMonitor_35_or73 | TLMonitor_35_or74;
  assign TLMonitor_35_or17 = TLMonitor_35_or35 | TLMonitor_35_or36;
  assign TLMonitor_35_or75 = stopEn33 | stopEn34;
  assign TLMonitor_35_or154 = stopEn36 | stopEn37;
  assign TLMonitor_35_or76 = stopEn35 | TLMonitor_35_or154;
  assign TLMonitor_35_or37 = TLMonitor_35_or75 | TLMonitor_35_or76;
  assign TLMonitor_35_or156 = stopEn39 | stopEn40;
  assign TLMonitor_35_or77 = stopEn38 | TLMonitor_35_or156;
  assign TLMonitor_35_or158 = stopEn42 | stopEn43;
  assign TLMonitor_35_or78 = stopEn41 | TLMonitor_35_or158;
  assign TLMonitor_35_or38 = TLMonitor_35_or77 | TLMonitor_35_or78;
  assign TLMonitor_35_or18 = TLMonitor_35_or37 | TLMonitor_35_or38;
  assign TLMonitor_35_or8 = TLMonitor_35_or17 | TLMonitor_35_or18;
  assign TLMonitor_35_or3 = TLMonitor_35_or7 | TLMonitor_35_or8;
  assign TLMonitor_35_or79 = stopEn44 | stopEn45;
  assign TLMonitor_35_or162 = stopEn47 | stopEn48;
  assign TLMonitor_35_or80 = stopEn46 | TLMonitor_35_or162;
  assign TLMonitor_35_or39 = TLMonitor_35_or79 | TLMonitor_35_or80;
  assign TLMonitor_35_or164 = stopEn50 | stopEn51;
  assign TLMonitor_35_or81 = stopEn49 | TLMonitor_35_or164;
  assign TLMonitor_35_or166 = stopEn53 | stopEn54;
  assign TLMonitor_35_or82 = stopEn52 | TLMonitor_35_or166;
  assign TLMonitor_35_or40 = TLMonitor_35_or81 | TLMonitor_35_or82;
  assign TLMonitor_35_or19 = TLMonitor_35_or39 | TLMonitor_35_or40;
  assign TLMonitor_35_or83 = stopEn55 | stopEn56;
  assign TLMonitor_35_or170 = stopEn58 | stopEn59;
  assign TLMonitor_35_or84 = stopEn57 | TLMonitor_35_or170;
  assign TLMonitor_35_or41 = TLMonitor_35_or83 | TLMonitor_35_or84;
  assign TLMonitor_35_or172 = stopEn61 | stopEn62;
  assign TLMonitor_35_or85 = stopEn60 | TLMonitor_35_or172;
  assign TLMonitor_35_or174 = stopEn64 | stopEn65;
  assign TLMonitor_35_or86 = stopEn63 | TLMonitor_35_or174;
  assign TLMonitor_35_or42 = TLMonitor_35_or85 | TLMonitor_35_or86;
  assign TLMonitor_35_or20 = TLMonitor_35_or41 | TLMonitor_35_or42;
  assign TLMonitor_35_or9 = TLMonitor_35_or19 | TLMonitor_35_or20;
  assign TLMonitor_35_or87 = stopEn66 | stopEn67;
  assign TLMonitor_35_or178 = stopEn69 | stopEn70;
  assign TLMonitor_35_or88 = stopEn68 | TLMonitor_35_or178;
  assign TLMonitor_35_or43 = TLMonitor_35_or87 | TLMonitor_35_or88;
  assign TLMonitor_35_or180 = stopEn72 | stopEn73;
  assign TLMonitor_35_or89 = stopEn71 | TLMonitor_35_or180;
  assign TLMonitor_35_or182 = stopEn75 | stopEn76;
  assign TLMonitor_35_or90 = stopEn74 | TLMonitor_35_or182;
  assign TLMonitor_35_or44 = TLMonitor_35_or89 | TLMonitor_35_or90;
  assign TLMonitor_35_or21 = TLMonitor_35_or43 | TLMonitor_35_or44;
  assign TLMonitor_35_or91 = stopEn77 | stopEn78;
  assign TLMonitor_35_or186 = stopEn80 | stopEn81;
  assign TLMonitor_35_or92 = stopEn79 | TLMonitor_35_or186;
  assign TLMonitor_35_or45 = TLMonitor_35_or91 | TLMonitor_35_or92;
  assign TLMonitor_35_or188 = stopEn83 | stopEn84;
  assign TLMonitor_35_or93 = stopEn82 | TLMonitor_35_or188;
  assign TLMonitor_35_or190 = stopEn86 | stopEn87;
  assign TLMonitor_35_or94 = stopEn85 | TLMonitor_35_or190;
  assign TLMonitor_35_or46 = TLMonitor_35_or93 | TLMonitor_35_or94;
  assign TLMonitor_35_or22 = TLMonitor_35_or45 | TLMonitor_35_or46;
  assign TLMonitor_35_or10 = TLMonitor_35_or21 | TLMonitor_35_or22;
  assign TLMonitor_35_or4 = TLMonitor_35_or9 | TLMonitor_35_or10;
  assign TLMonitor_35_or1 = TLMonitor_35_or3 | TLMonitor_35_or4;
  assign TLMonitor_35_or95 = stopEn88 | stopEn89;
  assign TLMonitor_35_or194 = stopEn91 | stopEn92;
  assign TLMonitor_35_or96 = stopEn90 | TLMonitor_35_or194;
  assign TLMonitor_35_or47 = TLMonitor_35_or95 | TLMonitor_35_or96;
  assign TLMonitor_35_or196 = stopEn94 | stopEn95;
  assign TLMonitor_35_or97 = stopEn93 | TLMonitor_35_or196;
  assign TLMonitor_35_or198 = stopEn97 | stopEn98;
  assign TLMonitor_35_or98 = stopEn96 | TLMonitor_35_or198;
  assign TLMonitor_35_or48 = TLMonitor_35_or97 | TLMonitor_35_or98;
  assign TLMonitor_35_or23 = TLMonitor_35_or47 | TLMonitor_35_or48;
  assign TLMonitor_35_or99 = stopEn99 | stopEn100;
  assign TLMonitor_35_or202 = stopEn102 | stopEn103;
  assign TLMonitor_35_or100 = stopEn101 | TLMonitor_35_or202;
  assign TLMonitor_35_or49 = TLMonitor_35_or99 | TLMonitor_35_or100;
  assign TLMonitor_35_or204 = stopEn105 | stopEn106;
  assign TLMonitor_35_or101 = stopEn104 | TLMonitor_35_or204;
  assign TLMonitor_35_or206 = stopEn108 | stopEn109;
  assign TLMonitor_35_or102 = stopEn107 | TLMonitor_35_or206;
  assign TLMonitor_35_or50 = TLMonitor_35_or101 | TLMonitor_35_or102;
  assign TLMonitor_35_or24 = TLMonitor_35_or49 | TLMonitor_35_or50;
  assign TLMonitor_35_or11 = TLMonitor_35_or23 | TLMonitor_35_or24;
  assign TLMonitor_35_or103 = stopEn110 | stopEn111;
  assign TLMonitor_35_or210 = stopEn113 | stopEn114;
  assign TLMonitor_35_or104 = stopEn112 | TLMonitor_35_or210;
  assign TLMonitor_35_or51 = TLMonitor_35_or103 | TLMonitor_35_or104;
  assign TLMonitor_35_or212 = stopEn116 | stopEn117;
  assign TLMonitor_35_or105 = stopEn115 | TLMonitor_35_or212;
  assign TLMonitor_35_or214 = stopEn119 | stopEn120;
  assign TLMonitor_35_or106 = stopEn118 | TLMonitor_35_or214;
  assign TLMonitor_35_or52 = TLMonitor_35_or105 | TLMonitor_35_or106;
  assign TLMonitor_35_or25 = TLMonitor_35_or51 | TLMonitor_35_or52;
  assign TLMonitor_35_or107 = stopEn121 | stopEn122;
  assign TLMonitor_35_or218 = stopEn124 | stopEn125;
  assign TLMonitor_35_or108 = stopEn123 | TLMonitor_35_or218;
  assign TLMonitor_35_or53 = TLMonitor_35_or107 | TLMonitor_35_or108;
  assign TLMonitor_35_or220 = stopEn127 | stopEn128;
  assign TLMonitor_35_or109 = stopEn126 | TLMonitor_35_or220;
  assign TLMonitor_35_or222 = stopEn130 | stopEn131;
  assign TLMonitor_35_or110 = stopEn129 | TLMonitor_35_or222;
  assign TLMonitor_35_or54 = TLMonitor_35_or109 | TLMonitor_35_or110;
  assign TLMonitor_35_or26 = TLMonitor_35_or53 | TLMonitor_35_or54;
  assign TLMonitor_35_or12 = TLMonitor_35_or25 | TLMonitor_35_or26;
  assign TLMonitor_35_or5 = TLMonitor_35_or11 | TLMonitor_35_or12;
  assign TLMonitor_35_or111 = stopEn132 | stopEn133;
  assign TLMonitor_35_or226 = stopEn135 | stopEn136;
  assign TLMonitor_35_or112 = stopEn134 | TLMonitor_35_or226;
  assign TLMonitor_35_or55 = TLMonitor_35_or111 | TLMonitor_35_or112;
  assign TLMonitor_35_or228 = stopEn138 | stopEn139;
  assign TLMonitor_35_or113 = stopEn137 | TLMonitor_35_or228;
  assign TLMonitor_35_or230 = stopEn141 | stopEn142;
  assign TLMonitor_35_or114 = stopEn140 | TLMonitor_35_or230;
  assign TLMonitor_35_or56 = TLMonitor_35_or113 | TLMonitor_35_or114;
  assign TLMonitor_35_or27 = TLMonitor_35_or55 | TLMonitor_35_or56;
  assign TLMonitor_35_or115 = stopEn143 | stopEn144;
  assign TLMonitor_35_or234 = stopEn146 | stopEn147;
  assign TLMonitor_35_or116 = stopEn145 | TLMonitor_35_or234;
  assign TLMonitor_35_or57 = TLMonitor_35_or115 | TLMonitor_35_or116;
  assign TLMonitor_35_or236 = stopEn149 | stopEn150;
  assign TLMonitor_35_or117 = stopEn148 | TLMonitor_35_or236;
  assign TLMonitor_35_or238 = stopEn152 | stopEn153;
  assign TLMonitor_35_or118 = stopEn151 | TLMonitor_35_or238;
  assign TLMonitor_35_or58 = TLMonitor_35_or117 | TLMonitor_35_or118;
  assign TLMonitor_35_or28 = TLMonitor_35_or57 | TLMonitor_35_or58;
  assign TLMonitor_35_or13 = TLMonitor_35_or27 | TLMonitor_35_or28;
  assign TLMonitor_35_or119 = stopEn154 | stopEn155;
  assign TLMonitor_35_or242 = stopEn157 | stopEn158;
  assign TLMonitor_35_or120 = stopEn156 | TLMonitor_35_or242;
  assign TLMonitor_35_or59 = TLMonitor_35_or119 | TLMonitor_35_or120;
  assign TLMonitor_35_or244 = stopEn160 | stopEn161;
  assign TLMonitor_35_or121 = stopEn159 | TLMonitor_35_or244;
  assign TLMonitor_35_or246 = stopEn163 | stopEn164;
  assign TLMonitor_35_or122 = stopEn162 | TLMonitor_35_or246;
  assign TLMonitor_35_or60 = TLMonitor_35_or121 | TLMonitor_35_or122;
  assign TLMonitor_35_or29 = TLMonitor_35_or59 | TLMonitor_35_or60;
  assign TLMonitor_35_or123 = stopEn165 | stopEn166;
  assign TLMonitor_35_or250 = stopEn168 | stopEn169;
  assign TLMonitor_35_or124 = stopEn167 | TLMonitor_35_or250;
  assign TLMonitor_35_or61 = TLMonitor_35_or123 | TLMonitor_35_or124;
  assign TLMonitor_35_or252 = stopEn171 | stopEn172;
  assign TLMonitor_35_or125 = stopEn170 | TLMonitor_35_or252;
  assign TLMonitor_35_or254 = stopEn174 | stopEn175;
  assign TLMonitor_35_or126 = stopEn173 | TLMonitor_35_or254;
  assign TLMonitor_35_or62 = TLMonitor_35_or125 | TLMonitor_35_or126;
  assign TLMonitor_35_or30 = TLMonitor_35_or61 | TLMonitor_35_or62;
  assign TLMonitor_35_or14 = TLMonitor_35_or29 | TLMonitor_35_or30;
  assign TLMonitor_35_or6 = TLMonitor_35_or13 | TLMonitor_35_or14;
  assign TLMonitor_35_or2 = TLMonitor_35_or5 | TLMonitor_35_or6;
  assign TLMonitor_35_or0 = TLMonitor_35_or1 | TLMonitor_35_or2;
  assign metaAssert = TLMonitor_35_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1575 = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1586 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1587 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1588 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1589 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1590 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1623 = _RAND_6[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1634 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1635 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1636 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1637 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_1638 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1639 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_1677 = _RAND_13[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_1688 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_1689 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1690 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_1691 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_1692 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_1725 = _RAND_19[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_1736 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_1737 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_1738 = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_1739 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_1740 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  inflight = _RAND_25[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  inflight_opcodes = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  inflight_sizes = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_1774 = _RAND_28[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_1792 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_1935 = _RAND_30[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_1944 = _RAND_31[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  TLMonitor_35_metaAssert = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_1575 <= 9'h0;
    end else if (reset) begin
      _T_1575 <= 9'h0;
    end else if (_T_1566) begin
      if (_T_1578) begin
        if (~io_in_a_bits_opcode[2]) begin
          _T_1575 <= _T_1571;
        end else begin
          _T_1575 <= 9'h0;
        end
      end else begin
        _T_1575 <= _T_1577;
      end
    end
    if (metaReset) begin
      _T_1586 <= 3'h0;
    end else if (_T_1614) begin
      _T_1586 <= io_in_a_bits_opcode;
    end
    if (metaReset) begin
      _T_1587 <= 3'h0;
    end else if (_T_1614) begin
      _T_1587 <= io_in_a_bits_param;
    end
    if (metaReset) begin
      _T_1588 <= 4'h0;
    end else if (_T_1614) begin
      _T_1588 <= io_in_a_bits_size;
    end
    if (metaReset) begin
      _T_1589 <= 1'h0;
    end else if (_T_1614) begin
      _T_1589 <= io_in_a_bits_source;
    end
    if (metaReset) begin
      _T_1590 <= 32'h0;
    end else if (_T_1614) begin
      _T_1590 <= io_in_a_bits_address;
    end
    if (metaReset) begin
      _T_1623 <= 9'h0;
    end else if (reset) begin
      _T_1623 <= 9'h0;
    end else if (_T_1615) begin
      if (_T_1626) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1623 <= _T_1620;
        end else begin
          _T_1623 <= 9'h0;
        end
      end else begin
        _T_1623 <= _T_1625;
      end
    end
    if (metaReset) begin
      _T_1634 <= 3'h0;
    end else if (_T_1667) begin
      _T_1634 <= io_in_d_bits_opcode;
    end
    if (metaReset) begin
      _T_1635 <= 2'h0;
    end else if (_T_1667) begin
      _T_1635 <= io_in_d_bits_param;
    end
    if (metaReset) begin
      _T_1636 <= 4'h0;
    end else if (_T_1667) begin
      _T_1636 <= io_in_d_bits_size;
    end
    if (metaReset) begin
      _T_1637 <= 1'h0;
    end else if (_T_1667) begin
      _T_1637 <= io_in_d_bits_source;
    end
    if (metaReset) begin
      _T_1638 <= 2'h0;
    end else if (_T_1667) begin
      _T_1638 <= io_in_d_bits_sink;
    end
    if (metaReset) begin
      _T_1639 <= 1'h0;
    end else if (_T_1667) begin
      _T_1639 <= io_in_d_bits_denied;
    end
    if (metaReset) begin
      _T_1677 <= 9'h0;
    end else if (reset) begin
      _T_1677 <= 9'h0;
    end else if (_T_1668) begin
      if (_T_1680) begin
        _T_1677 <= 9'h0;
      end else begin
        _T_1677 <= _T_1679;
      end
    end
    if (metaReset) begin
      _T_1688 <= 3'h0;
    end else if (_T_1716) begin
      _T_1688 <= io_in_b_bits_opcode;
    end
    if (metaReset) begin
      _T_1689 <= 2'h0;
    end else if (_T_1716) begin
      _T_1689 <= io_in_b_bits_param;
    end
    if (metaReset) begin
      _T_1690 <= 4'h0;
    end else if (_T_1716) begin
      _T_1690 <= io_in_b_bits_size;
    end
    if (metaReset) begin
      _T_1691 <= 1'h0;
    end else if (_T_1716) begin
      _T_1691 <= io_in_b_bits_source;
    end
    if (metaReset) begin
      _T_1692 <= 32'h0;
    end else if (_T_1716) begin
      _T_1692 <= io_in_b_bits_address;
    end
    if (metaReset) begin
      _T_1725 <= 9'h0;
    end else if (reset) begin
      _T_1725 <= 9'h0;
    end else if (_T_1717) begin
      if (_T_1728) begin
        if (io_in_c_bits_opcode[0]) begin
          _T_1725 <= _T_1722;
        end else begin
          _T_1725 <= 9'h0;
        end
      end else begin
        _T_1725 <= _T_1727;
      end
    end
    if (metaReset) begin
      _T_1736 <= 3'h0;
    end else if (_T_1764) begin
      _T_1736 <= io_in_c_bits_opcode;
    end
    if (metaReset) begin
      _T_1737 <= 3'h0;
    end else if (_T_1764) begin
      _T_1737 <= io_in_c_bits_param;
    end
    if (metaReset) begin
      _T_1738 <= 4'h0;
    end else if (_T_1764) begin
      _T_1738 <= io_in_c_bits_size;
    end
    if (metaReset) begin
      _T_1739 <= 1'h0;
    end else if (_T_1764) begin
      _T_1739 <= io_in_c_bits_source;
    end
    if (metaReset) begin
      _T_1740 <= 32'h0;
    end else if (_T_1764) begin
      _T_1740 <= io_in_c_bits_address;
    end
    if (metaReset) begin
      inflight <= 2'h0;
    end else if (reset) begin
      inflight <= 2'h0;
    end else begin
      inflight <= _T_1913;
    end
    if (metaReset) begin
      inflight_opcodes <= 8'h0;
    end else if (reset) begin
      inflight_opcodes <= 8'h0;
    end else begin
      inflight_opcodes <= _T_1916;
    end
    if (metaReset) begin
      inflight_sizes <= 16'h0;
    end else if (reset) begin
      inflight_sizes <= 16'h0;
    end else begin
      inflight_sizes <= _T_1919;
    end
    if (metaReset) begin
      _T_1774 <= 9'h0;
    end else if (reset) begin
      _T_1774 <= 9'h0;
    end else if (_T_1566) begin
      if (a_first) begin
        if (~io_in_a_bits_opcode[2]) begin
          _T_1774 <= _T_1571;
        end else begin
          _T_1774 <= 9'h0;
        end
      end else begin
        _T_1774 <= _T_1776;
      end
    end
    if (metaReset) begin
      _T_1792 <= 9'h0;
    end else if (reset) begin
      _T_1792 <= 9'h0;
    end else if (_T_1615) begin
      if (d_first) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1792 <= _T_1620;
        end else begin
          _T_1792 <= 9'h0;
        end
      end else begin
        _T_1792 <= _T_1794;
      end
    end
    if (metaReset) begin
      _T_1935 <= 4'h0;
    end else if (reset) begin
      _T_1935 <= 4'h0;
    end else begin
      _T_1935 <= _T_1983;
    end
    if (metaReset) begin
      _T_1944 <= 9'h0;
    end else if (reset) begin
      _T_1944 <= 9'h0;
    end else if (_T_1615) begin
      if (_T_1947) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1944 <= _T_1620;
        end else begin
          _T_1944 <= 9'h0;
        end
      end else begin
        _T_1944 <= _T_1946;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & ~_T_128) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & ~_T_128) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & ~_T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & ~_T_151) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & ~_T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & ~_T_154) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & ~_T_158) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & ~_T_158) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & ~_T_161) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & ~_T_161) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & ~_T_165) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & ~_T_165) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & ~_T_170) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & ~_T_170) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & ~_T_128) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & ~_T_128) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & ~_T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & ~_T_151) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & ~_T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & ~_T_154) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & ~_T_158) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & ~_T_158) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & ~_T_161) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & ~_T_161) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & ~_T_165) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & ~_T_165) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & ~_T_247) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & ~_T_247) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & ~_T_170) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & ~_T_170) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & ~_T_321) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type which is unexpected using diplomatic parameters\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & ~_T_321) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & ~_T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & ~_T_154) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & ~_T_161) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & ~_T_161) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & ~_T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & ~_T_331) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & ~_T_335) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & ~_T_335) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_411) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_154) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_161) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_161) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_331) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_335) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_335) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_135 & ~_T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_135 & ~_T_411) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_135 & ~_T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_135 & ~_T_154) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_135 & ~_T_161) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_135 & ~_T_161) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_135 & ~_T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_135 & ~_T_331) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_135 & ~_T_513) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_135 & ~_T_513) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & ~_T_563) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & ~_T_563) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & ~_T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & ~_T_154) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & ~_T_161) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & ~_T_161) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & ~_T_573) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & ~_T_573) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & ~_T_335) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & ~_T_335) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & ~_T_563) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & ~_T_563) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & ~_T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & ~_T_154) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & ~_T_161) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & ~_T_161) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & ~_T_637) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & ~_T_637) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & ~_T_335) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & ~_T_335) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & ~_T_703) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & ~_T_703) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & ~_T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & ~_T_154) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & ~_T_161) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & ~_T_161) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & ~_T_713) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid opcode param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & ~_T_713) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & ~_T_335) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & ~_T_335) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~_T_725) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~_T_725) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & ~_T_734) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & ~_T_734) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & ~_T_738) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & ~_T_738) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & ~_T_742) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & ~_T_742) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & ~_T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & ~_T_746) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & ~_T_750) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & ~_T_750) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & ~_T_734) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & ~_T_734) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & ~_T_738) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & ~_T_738) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & ~_T_765) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & ~_T_765) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & ~_T_769) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & ~_T_769) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & ~_T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & ~_T_746) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_734) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_734) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_738) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_738) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_765) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_765) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_769) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_769) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_802) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_802) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & ~_T_734) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & ~_T_734) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & ~_T_742) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & ~_T_742) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & ~_T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & ~_T_746) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & ~_T_734) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & ~_T_734) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & ~_T_742) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & ~_T_742) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & ~_T_802) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & ~_T_802) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_217 & ~_T_734) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_217 & ~_T_734) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_217 & ~_T_742) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_217 & ~_T_742) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_217 & ~_T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_217 & ~_T_746) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & ~_T_863) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & ~_T_863) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & ~_T_1027) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type which is unexpected using diplomatic parameters (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & ~_T_1027) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & ~_T_1030) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & ~_T_1030) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & ~_T_1036) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & ~_T_1036) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & ~_T_1040) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & ~_T_1040) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & ~_T_1044) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & ~_T_1044) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & ~_T_1048) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & ~_T_1048) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_237 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type which is unexpected using diplomatic parameters (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_237 & ~reset) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_237 & ~_T_1030) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_237 & ~_T_1030) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_237 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_237 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_237 & ~_T_1036) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_237 & ~_T_1036) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_237 & ~_T_1077) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_237 & ~_T_1077) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_237 & ~_T_1044) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_237 & ~_T_1044) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_237 & ~_T_1048) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_237 & ~_T_1048) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type which is unexpected using diplomatic parameters (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~reset) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~_T_1030) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~_T_1030) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~_T_1036) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~_T_1036) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~_T_1077) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~_T_1077) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~_T_1044) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~_T_1044) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_263 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_263 & ~reset) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_263 & ~_T_1030) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_263 & ~_T_1030) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_263 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_263 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_263 & ~_T_1036) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_263 & ~_T_1036) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_263 & ~_T_1077) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_263 & ~_T_1077) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_263 & ~_T_1153) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_263 & ~_T_1153) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by master (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & ~reset) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & ~_T_1030) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & ~_T_1030) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & ~_T_1036) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & ~_T_1036) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & ~_T_1044) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & ~_T_1044) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~reset) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1030) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1030) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1036) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1036) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1044) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1044) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & ~reset) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & ~_T_1030) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & ~_T_1030) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & ~_T_1036) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & ~_T_1036) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & ~_T_1044) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & ~_T_1044) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & ~_T_1048) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & ~_T_1048) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_307 & ~_T_1332) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_307 & ~_T_1332) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_307 & ~_T_1335) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_307 & ~_T_1335) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_307 & ~_T_1339) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_307 & ~_T_1339) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_307 & ~_T_1342) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_307 & ~_T_1342) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_307 & ~_T_1346) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_307 & ~_T_1346) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1332) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1332) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1335) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1335) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1339) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1339) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1342) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1342) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1346) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1346) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & ~_T_1400) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & ~_T_1400) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & ~_T_1423) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & ~_T_1423) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & ~_T_1335) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & ~_T_1335) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & ~_T_1339) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & ~_T_1339) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & ~_T_1342) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & ~_T_1342) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & ~_T_1437) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & ~_T_1437) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_339 & ~_T_1400) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_339 & ~_T_1400) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_339 & ~_T_1423) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_339 & ~_T_1423) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_339 & ~_T_1335) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_339 & ~_T_1335) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_339 & ~_T_1339) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_339 & ~_T_1339) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_339 & ~_T_1342) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_339 & ~_T_1342) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_339 & ~_T_1437) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_339 & ~_T_1437) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_351 & ~_T_1332) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_351 & ~_T_1332) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_351 & ~_T_1335) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_351 & ~_T_1335) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_351 & ~_T_1342) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_351 & ~_T_1342) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_351 & ~_T_1524) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_351 & ~_T_1524) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_359 & ~_T_1332) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_359 & ~_T_1332) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_359 & ~_T_1335) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_359 & ~_T_1335) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_359 & ~_T_1342) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_359 & ~_T_1342) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_359 & ~_T_1524) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_359 & ~_T_1524) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & ~_T_1332) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_367 & ~_T_1332) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & ~_T_1335) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_367 & ~_T_1335) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & ~_T_1342) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_367 & ~_T_1342) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & ~_T_1524) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_367 & ~_T_1524) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1592 & ~_T_1595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1592 & ~_T_1595) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1592 & ~_T_1599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1592 & ~_T_1599) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1592 & ~_T_1603) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1592 & ~_T_1603) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1592 & ~_T_1607) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1592 & ~_T_1607) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1592 & ~_T_1611) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1592 & ~_T_1611) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1641 & ~_T_1644) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1641 & ~_T_1644) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1641 & ~_T_1648) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1641 & ~_T_1648) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1641 & ~_T_1652) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1641 & ~_T_1652) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1641 & ~_T_1656) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1641 & ~_T_1656) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1641 & ~_T_1660) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1641 & ~_T_1660) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1641 & ~_T_1664) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1641 & ~_T_1664) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1694 & ~_T_1697) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1694 & ~_T_1697) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1694 & ~_T_1701) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1694 & ~_T_1701) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1694 & ~_T_1705) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1694 & ~_T_1705) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1694 & ~_T_1709) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1694 & ~_T_1709) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1694 & ~_T_1713) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1694 & ~_T_1713) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1742 & ~_T_1745) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1742 & ~_T_1745) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1742 & ~_T_1749) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1742 & ~_T_1749) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1742 & ~_T_1753) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1742 & ~_T_1753) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1742 & ~_T_1757) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1742 & ~_T_1757) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1742 & ~_T_1761) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1742 & ~_T_1761) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1821 & ~_T_1836) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1821 & ~_T_1836) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1860 & ~_T_1870) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1860 & ~_T_1870) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1860 & ~_T_1883) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1860 & ~_T_1883) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1860 & ~_T_1890) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1860 & ~_T_1890) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1898 & ~_T_1902) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1898 & ~_T_1902) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1909) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1909) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1962 & ~_T_1968) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at HellaCache.scala:256:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1962 & ~_T_1968) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1971 & ~_T_1979) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at HellaCache.scala:256:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1971 & ~_T_1979) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    if (metaReset) begin
      TLMonitor_35_metaAssert <= 1'h0;
    end else begin
      TLMonitor_35_metaAssert <= TLMonitor_35_metaAssert | TLMonitor_35_or0;
    end
  end
endmodule
module TLMonitor_36(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [31:0] io_in_a_bits_address,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [3:0]  io_in_d_bits_size,
  input  [1:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [31:0] _T_10; // @[Edges.scala 22:16]
  wire  _T_11; // @[Edges.scala 22:24]
  wire [32:0] _T_79; // @[Parameters.scala 137:49]
  wire [31:0] _T_105; // @[Parameters.scala 137:31]
  wire [32:0] _T_106; // @[Parameters.scala 137:49]
  wire  _T_140; // @[Monitor.scala 44:11]
  wire [31:0] _T_238; // @[Parameters.scala 137:31]
  wire [32:0] _T_239; // @[Parameters.scala 137:49]
  wire [32:0] _T_241; // @[Parameters.scala 137:52]
  wire  _T_242; // @[Parameters.scala 137:67]
  wire [32:0] _T_251; // @[Parameters.scala 137:52]
  wire  _T_252; // @[Parameters.scala 137:67]
  wire [31:0] _T_253; // @[Parameters.scala 137:31]
  wire [32:0] _T_254; // @[Parameters.scala 137:49]
  wire [32:0] _T_256; // @[Parameters.scala 137:52]
  wire  _T_257; // @[Parameters.scala 137:67]
  wire [31:0] _T_258; // @[Parameters.scala 137:31]
  wire [32:0] _T_259; // @[Parameters.scala 137:49]
  wire [32:0] _T_261; // @[Parameters.scala 137:52]
  wire  _T_262; // @[Parameters.scala 137:67]
  wire [31:0] _T_263; // @[Parameters.scala 137:31]
  wire [32:0] _T_264; // @[Parameters.scala 137:49]
  wire [32:0] _T_266; // @[Parameters.scala 137:52]
  wire  _T_267; // @[Parameters.scala 137:67]
  wire [31:0] _T_268; // @[Parameters.scala 137:31]
  wire [32:0] _T_269; // @[Parameters.scala 137:49]
  wire [32:0] _T_271; // @[Parameters.scala 137:52]
  wire  _T_272; // @[Parameters.scala 137:67]
  wire [32:0] _T_276; // @[Parameters.scala 137:52]
  wire  _T_277; // @[Parameters.scala 137:67]
  wire  _T_278; // @[Parameters.scala 602:42]
  wire  _T_279; // @[Parameters.scala 602:42]
  wire  _T_280; // @[Parameters.scala 602:42]
  wire  _T_281; // @[Parameters.scala 602:42]
  wire  _T_282; // @[Parameters.scala 602:42]
  wire  _T_285; // @[Parameters.scala 603:30]
  wire  _T_288; // @[Monitor.scala 44:11]
  wire  _T_680; // @[Bundles.scala 44:24]
  wire  _T_682; // @[Monitor.scala 51:11]
  wire  _T_687; // @[Monitor.scala 310:25]
  wire  _T_691; // @[Monitor.scala 312:27]
  wire  _T_693; // @[Monitor.scala 51:11]
  wire  _T_695; // @[Monitor.scala 313:28]
  wire  _T_697; // @[Monitor.scala 51:11]
  wire  _T_701; // @[Monitor.scala 51:11]
  wire  _T_705; // @[Monitor.scala 51:11]
  wire  _T_707; // @[Monitor.scala 318:25]
  wire  _T_718; // @[Bundles.scala 104:26]
  wire  _T_720; // @[Monitor.scala 51:11]
  wire  _T_722; // @[Monitor.scala 323:28]
  wire  _T_724; // @[Monitor.scala 51:11]
  wire  _T_735; // @[Monitor.scala 328:25]
  wire  _T_755; // @[Monitor.scala 334:30]
  wire  _T_757; // @[Monitor.scala 51:11]
  wire  _T_764; // @[Monitor.scala 338:25]
  wire  _T_781; // @[Monitor.scala 346:25]
  wire  _T_799; // @[Monitor.scala 354:25]
  wire  _T_831; // @[Decoupled.scala 40:37]
  reg [8:0] _T_840; // @[Edges.scala 230:27]
  reg [31:0] _RAND_0;
  wire [8:0] _T_842; // @[Edges.scala 231:28]
  wire  _T_843; // @[Edges.scala 232:25]
  reg [31:0] _T_855; // @[Monitor.scala 388:22]
  reg [31:0] _RAND_1;
  wire  _T_857; // @[Monitor.scala 389:19]
  wire  _T_874; // @[Monitor.scala 394:32]
  wire  _T_876; // @[Monitor.scala 44:11]
  wire  _T_879; // @[Monitor.scala 396:20]
  wire [26:0] _T_882; // @[package.scala 212:77]
  wire [8:0] _T_885; // @[Edges.scala 221:59]
  reg [8:0] _T_888; // @[Edges.scala 230:27]
  reg [31:0] _RAND_2;
  wire [8:0] _T_890; // @[Edges.scala 231:28]
  wire  _T_891; // @[Edges.scala 232:25]
  reg [2:0] _T_899; // @[Monitor.scala 535:22]
  reg [31:0] _RAND_3;
  reg [1:0] _T_900; // @[Monitor.scala 536:22]
  reg [31:0] _RAND_4;
  reg [3:0] _T_901; // @[Monitor.scala 537:22]
  reg [31:0] _RAND_5;
  reg [1:0] _T_903; // @[Monitor.scala 539:22]
  reg [31:0] _RAND_6;
  reg  _T_904; // @[Monitor.scala 540:22]
  reg [31:0] _RAND_7;
  wire  _T_906; // @[Monitor.scala 541:19]
  wire  _T_907; // @[Monitor.scala 542:29]
  wire  _T_909; // @[Monitor.scala 51:11]
  wire  _T_911; // @[Monitor.scala 543:29]
  wire  _T_913; // @[Monitor.scala 51:11]
  wire  _T_915; // @[Monitor.scala 544:29]
  wire  _T_917; // @[Monitor.scala 51:11]
  wire  _T_923; // @[Monitor.scala 546:29]
  wire  _T_925; // @[Monitor.scala 51:11]
  wire  _T_927; // @[Monitor.scala 547:29]
  wire  _T_929; // @[Monitor.scala 51:11]
  wire  _T_932; // @[Monitor.scala 549:20]
  reg  inflight; // @[Monitor.scala 611:27]
  reg [31:0] _RAND_8;
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [31:0] _RAND_9;
  reg [7:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [31:0] _RAND_10;
  reg [8:0] _T_942; // @[Edges.scala 230:27]
  reg [31:0] _RAND_11;
  wire [8:0] _T_944; // @[Edges.scala 231:28]
  wire  a_first; // @[Edges.scala 232:25]
  reg [8:0] _T_960; // @[Edges.scala 230:27]
  reg [31:0] _RAND_12;
  wire [8:0] _T_962; // @[Edges.scala 231:28]
  wire  d_first; // @[Edges.scala 232:25]
  wire [15:0] _T_975; // @[Monitor.scala 609:57]
  wire [15:0] _GEN_56; // @[Monitor.scala 632:97]
  wire [15:0] _T_976; // @[Monitor.scala 632:97]
  wire [15:0] _T_977; // @[Monitor.scala 632:152]
  wire [15:0] _T_983; // @[Monitor.scala 609:57]
  wire [15:0] _GEN_58; // @[Monitor.scala 636:91]
  wire [15:0] _T_984; // @[Monitor.scala 636:91]
  wire [15:0] _T_985; // @[Monitor.scala 636:144]
  wire  _T_989; // @[Monitor.scala 646:27]
  wire [3:0] a_opcodes_set_interm; // @[Monitor.scala 646:72]
  wire [18:0] _T_997; // @[Monitor.scala 650:47]
  wire [4:0] a_sizes_set_interm; // @[Monitor.scala 646:72]
  wire [19:0] _T_999; // @[Monitor.scala 651:43]
  wire  _T_1004; // @[Monitor.scala 44:11]
  wire [1:0] _GEN_15; // @[Monitor.scala 646:72]
  wire [18:0] _GEN_18; // @[Monitor.scala 646:72]
  wire [19:0] _GEN_19; // @[Monitor.scala 646:72]
  wire  _T_1008; // @[Monitor.scala 663:27]
  wire  _T_1011; // @[Monitor.scala 663:72]
  wire [30:0] _T_1018; // @[Monitor.scala 665:76]
  wire [30:0] _T_1024; // @[Monitor.scala 666:72]
  wire [1:0] _GEN_20; // @[Monitor.scala 663:91]
  wire [30:0] _GEN_21; // @[Monitor.scala 663:91]
  wire [30:0] _GEN_22; // @[Monitor.scala 663:91]
  wire  _T_1033; // @[Monitor.scala 669:142]
  wire  _T_1034; // @[Monitor.scala 669:119]
  wire  _T_1035; // @[Monitor.scala 669:166]
  wire  _T_1036; // @[Monitor.scala 669:49]
  wire  _T_1038; // @[Monitor.scala 51:11]
  wire [3:0] a_opcode_lookup; // @[Monitor.scala 632:21]
  wire [2:0] _GEN_25; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_26; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_27; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_28; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_29; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_30; // @[Monitor.scala 670:37]
  wire  _T_1041; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_37; // @[Monitor.scala 670:96]
  wire [2:0] _GEN_38; // @[Monitor.scala 670:96]
  wire  _T_1043; // @[Monitor.scala 670:96]
  wire  _T_1044; // @[Monitor.scala 670:71]
  wire  _T_1047; // @[Monitor.scala 671:99]
  wire  _T_1048; // @[Monitor.scala 671:34]
  wire  _T_1049; // @[Monitor.scala 671:15]
  wire  _T_1051; // @[Monitor.scala 51:11]
  wire [7:0] a_size_lookup; // @[Monitor.scala 636:19]
  wire [7:0] _GEN_60; // @[Monitor.scala 673:34]
  wire  _T_1053; // @[Monitor.scala 673:34]
  wire  _T_1056; // @[Monitor.scala 673:53]
  wire  _T_1058; // @[Monitor.scala 51:11]
  wire  _T_1061; // @[Monitor.scala 675:36]
  wire  _T_1062; // @[Monitor.scala 675:47]
  wire  _T_1066; // @[Monitor.scala 675:116]
  wire  _T_1070; // @[Monitor.scala 51:11]
  wire  a_set; // @[Monitor.scala 647:13]
  wire  d_clr; // @[Monitor.scala 664:13]
  wire  _T_1072; // @[Monitor.scala 680:20]
  wire  _T_1073; // @[Monitor.scala 680:40]
  wire  _T_1075; // @[Monitor.scala 680:30]
  wire  _T_1077; // @[Monitor.scala 51:11]
  wire  _T_1079; // @[Monitor.scala 683:27]
  wire  _T_1081; // @[Monitor.scala 683:36]
  wire [3:0] a_opcodes_set; // @[Monitor.scala 650:21]
  wire [3:0] _T_1082; // @[Monitor.scala 684:43]
  wire [3:0] d_opcodes_clr; // @[Monitor.scala 665:21]
  wire [3:0] _T_1084; // @[Monitor.scala 684:60]
  wire [7:0] a_sizes_set; // @[Monitor.scala 651:19]
  wire [7:0] _T_1085; // @[Monitor.scala 685:39]
  wire [7:0] d_sizes_clr; // @[Monitor.scala 666:19]
  wire [7:0] _T_1087; // @[Monitor.scala 685:54]
  wire  _GEN_61; // @[Monitor.scala 51:11]
  wire  _GEN_69; // @[Monitor.scala 51:11]
  wire  _GEN_77; // @[Monitor.scala 51:11]
  wire  _GEN_85; // @[Monitor.scala 51:11]
  wire  _GEN_89; // @[Monitor.scala 51:11]
  wire  _GEN_93; // @[Monitor.scala 51:11]
  wire [29:0] TLMonitor_36_covSum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  stopEn4;
  wire  stopEn5;
  wire  stopEn6;
  wire  stopEn7;
  wire  stopEn8;
  wire  stopEn9;
  wire  stopEn10;
  wire  stopEn11;
  wire  stopEn12;
  wire  stopEn13;
  wire  stopEn14;
  wire  stopEn15;
  wire  stopEn16;
  wire  stopEn17;
  wire  stopEn18;
  wire  stopEn19;
  wire  stopEn20;
  wire  stopEn21;
  wire  stopEn22;
  wire  stopEn23;
  wire  stopEn24;
  wire  stopEn25;
  wire  stopEn26;
  wire  stopEn27;
  wire  stopEn28;
  wire  stopEn29;
  wire  stopEn30;
  wire  stopEn31;
  wire  stopEn32;
  wire  TLMonitor_36_or15;
  wire  TLMonitor_36_or16;
  wire  TLMonitor_36_or7;
  wire  TLMonitor_36_or17;
  wire  TLMonitor_36_or18;
  wire  TLMonitor_36_or8;
  wire  TLMonitor_36_or3;
  wire  TLMonitor_36_or19;
  wire  TLMonitor_36_or20;
  wire  TLMonitor_36_or9;
  wire  TLMonitor_36_or21;
  wire  TLMonitor_36_or22;
  wire  TLMonitor_36_or10;
  wire  TLMonitor_36_or4;
  wire  TLMonitor_36_or1;
  wire  TLMonitor_36_or23;
  wire  TLMonitor_36_or24;
  wire  TLMonitor_36_or11;
  wire  TLMonitor_36_or25;
  wire  TLMonitor_36_or26;
  wire  TLMonitor_36_or12;
  wire  TLMonitor_36_or5;
  wire  TLMonitor_36_or27;
  wire  TLMonitor_36_or28;
  wire  TLMonitor_36_or13;
  wire  TLMonitor_36_or29;
  wire  TLMonitor_36_or62;
  wire  TLMonitor_36_or30;
  wire  TLMonitor_36_or14;
  wire  TLMonitor_36_or6;
  wire  TLMonitor_36_or2;
  wire  TLMonitor_36_or0;
  reg  TLMonitor_36_metaAssert;
  reg [31:0] _RAND_13;
  assign _T_10 = io_in_a_bits_address & 32'h3f; // @[Edges.scala 22:16]
  assign _T_11 = _T_10 == 32'h0; // @[Edges.scala 22:24]
  assign _T_79 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49]
  assign _T_105 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  assign _T_106 = {1'b0,$signed(_T_105)}; // @[Parameters.scala 137:49]
  assign _T_140 = _T_11 | reset; // @[Monitor.scala 44:11]
  assign _T_238 = io_in_a_bits_address ^ 32'h2000; // @[Parameters.scala 137:31]
  assign _T_239 = {1'b0,$signed(_T_238)}; // @[Parameters.scala 137:49]
  assign _T_241 = $signed(_T_239) & 33'shca012000; // @[Parameters.scala 137:52]
  assign _T_242 = $signed(_T_241) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_251 = $signed(_T_79) & 33'shca012000; // @[Parameters.scala 137:52]
  assign _T_252 = $signed(_T_251) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_253 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31]
  assign _T_254 = {1'b0,$signed(_T_253)}; // @[Parameters.scala 137:49]
  assign _T_256 = $signed(_T_254) & 33'shca010000; // @[Parameters.scala 137:52]
  assign _T_257 = $signed(_T_256) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_258 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31]
  assign _T_259 = {1'b0,$signed(_T_258)}; // @[Parameters.scala 137:49]
  assign _T_261 = $signed(_T_259) & 33'shca010000; // @[Parameters.scala 137:52]
  assign _T_262 = $signed(_T_261) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_263 = io_in_a_bits_address ^ 32'h8000000; // @[Parameters.scala 137:31]
  assign _T_264 = {1'b0,$signed(_T_263)}; // @[Parameters.scala 137:49]
  assign _T_266 = $signed(_T_264) & 33'shc8000000; // @[Parameters.scala 137:52]
  assign _T_267 = $signed(_T_266) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_268 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  assign _T_269 = {1'b0,$signed(_T_268)}; // @[Parameters.scala 137:49]
  assign _T_271 = $signed(_T_269) & 33'shc0000000; // @[Parameters.scala 137:52]
  assign _T_272 = $signed(_T_271) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_276 = $signed(_T_106) & 33'shc0000000; // @[Parameters.scala 137:52]
  assign _T_277 = $signed(_T_276) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_278 = _T_252 | _T_257; // @[Parameters.scala 602:42]
  assign _T_279 = _T_278 | _T_262; // @[Parameters.scala 602:42]
  assign _T_280 = _T_279 | _T_267; // @[Parameters.scala 602:42]
  assign _T_281 = _T_280 | _T_272; // @[Parameters.scala 602:42]
  assign _T_282 = _T_281 | _T_277; // @[Parameters.scala 602:42]
  assign _T_285 = _T_242 | _T_282; // @[Parameters.scala 603:30]
  assign _T_288 = _T_285 | reset; // @[Monitor.scala 44:11]
  assign _T_680 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 44:24]
  assign _T_682 = _T_680 | reset; // @[Monitor.scala 51:11]
  assign _T_687 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  assign _T_691 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27]
  assign _T_693 = _T_691 | reset; // @[Monitor.scala 51:11]
  assign _T_695 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  assign _T_697 = _T_695 | reset; // @[Monitor.scala 51:11]
  assign _T_701 = ~io_in_d_bits_corrupt | reset; // @[Monitor.scala 51:11]
  assign _T_705 = ~io_in_d_bits_denied | reset; // @[Monitor.scala 51:11]
  assign _T_707 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  assign _T_718 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 104:26]
  assign _T_720 = _T_718 | reset; // @[Monitor.scala 51:11]
  assign _T_722 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  assign _T_724 = _T_722 | reset; // @[Monitor.scala 51:11]
  assign _T_735 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  assign _T_755 = ~io_in_d_bits_denied | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  assign _T_757 = _T_755 | reset; // @[Monitor.scala 51:11]
  assign _T_764 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  assign _T_781 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  assign _T_799 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  assign _T_831 = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  assign _T_842 = _T_840 - 9'h1; // @[Edges.scala 231:28]
  assign _T_843 = _T_840 == 9'h0; // @[Edges.scala 232:25]
  assign _T_857 = io_in_a_valid & ~_T_843; // @[Monitor.scala 389:19]
  assign _T_874 = io_in_a_bits_address == _T_855; // @[Monitor.scala 394:32]
  assign _T_876 = _T_874 | reset; // @[Monitor.scala 44:11]
  assign _T_879 = _T_831 & _T_843; // @[Monitor.scala 396:20]
  assign _T_882 = 27'hfff << io_in_d_bits_size; // @[package.scala 212:77]
  assign _T_885 = ~_T_882[11:3]; // @[Edges.scala 221:59]
  assign _T_890 = _T_888 - 9'h1; // @[Edges.scala 231:28]
  assign _T_891 = _T_888 == 9'h0; // @[Edges.scala 232:25]
  assign _T_906 = io_in_d_valid & ~_T_891; // @[Monitor.scala 541:19]
  assign _T_907 = io_in_d_bits_opcode == _T_899; // @[Monitor.scala 542:29]
  assign _T_909 = _T_907 | reset; // @[Monitor.scala 51:11]
  assign _T_911 = io_in_d_bits_param == _T_900; // @[Monitor.scala 543:29]
  assign _T_913 = _T_911 | reset; // @[Monitor.scala 51:11]
  assign _T_915 = io_in_d_bits_size == _T_901; // @[Monitor.scala 544:29]
  assign _T_917 = _T_915 | reset; // @[Monitor.scala 51:11]
  assign _T_923 = io_in_d_bits_sink == _T_903; // @[Monitor.scala 546:29]
  assign _T_925 = _T_923 | reset; // @[Monitor.scala 51:11]
  assign _T_927 = io_in_d_bits_denied == _T_904; // @[Monitor.scala 547:29]
  assign _T_929 = _T_927 | reset; // @[Monitor.scala 51:11]
  assign _T_932 = io_in_d_valid & _T_891; // @[Monitor.scala 549:20]
  assign _T_944 = _T_942 - 9'h1; // @[Edges.scala 231:28]
  assign a_first = _T_942 == 9'h0; // @[Edges.scala 232:25]
  assign _T_962 = _T_960 - 9'h1; // @[Edges.scala 231:28]
  assign d_first = _T_960 == 9'h0; // @[Edges.scala 232:25]
  assign _T_975 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  assign _GEN_56 = {{12'd0}, inflight_opcodes}; // @[Monitor.scala 632:97]
  assign _T_976 = _GEN_56 & _T_975; // @[Monitor.scala 632:97]
  assign _T_977 = {{1'd0}, _T_976[15:1]}; // @[Monitor.scala 632:152]
  assign _T_983 = 16'h100 - 16'h1; // @[Monitor.scala 609:57]
  assign _GEN_58 = {{8'd0}, inflight_sizes}; // @[Monitor.scala 636:91]
  assign _T_984 = _GEN_58 & _T_983; // @[Monitor.scala 636:91]
  assign _T_985 = {{1'd0}, _T_984[15:1]}; // @[Monitor.scala 636:144]
  assign _T_989 = _T_831 & a_first; // @[Monitor.scala 646:27]
  assign a_opcodes_set_interm = _T_989 ? 4'h9 : 4'h0; // @[Monitor.scala 646:72]
  assign _T_997 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 650:47]
  assign a_sizes_set_interm = _T_989 ? 5'hd : 5'h0; // @[Monitor.scala 646:72]
  assign _T_999 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 651:43]
  assign _T_1004 = ~inflight | reset; // @[Monitor.scala 44:11]
  assign _GEN_15 = _T_989 ? 2'h1 : 2'h0; // @[Monitor.scala 646:72]
  assign _GEN_18 = _T_989 ? _T_997 : 19'h0; // @[Monitor.scala 646:72]
  assign _GEN_19 = _T_989 ? _T_999 : 20'h0; // @[Monitor.scala 646:72]
  assign _T_1008 = io_in_d_valid & d_first; // @[Monitor.scala 663:27]
  assign _T_1011 = _T_1008 & ~_T_687; // @[Monitor.scala 663:72]
  assign _T_1018 = {{15'd0}, _T_975}; // @[Monitor.scala 665:76]
  assign _T_1024 = {{15'd0}, _T_983}; // @[Monitor.scala 666:72]
  assign _GEN_20 = _T_1011 ? 2'h1 : 2'h0; // @[Monitor.scala 663:91]
  assign _GEN_21 = _T_1011 ? _T_1018 : 31'h0; // @[Monitor.scala 663:91]
  assign _GEN_22 = _T_1011 ? _T_1024 : 31'h0; // @[Monitor.scala 663:91]
  assign _T_1033 = 4'h6 == io_in_d_bits_size; // @[Monitor.scala 669:142]
  assign _T_1034 = io_in_a_valid & _T_1033; // @[Monitor.scala 669:119]
  assign _T_1035 = _T_1034 & a_first; // @[Monitor.scala 669:166]
  assign _T_1036 = inflight | _T_1035; // @[Monitor.scala 669:49]
  assign _T_1038 = _T_1036 | reset; // @[Monitor.scala 51:11]
  assign a_opcode_lookup = _T_977[3:0]; // @[Monitor.scala 632:21]
  assign _GEN_25 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 670:37]
  assign _GEN_26 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_25; // @[Monitor.scala 670:37]
  assign _GEN_27 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_26; // @[Monitor.scala 670:37]
  assign _GEN_28 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_27; // @[Monitor.scala 670:37]
  assign _GEN_29 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_28; // @[Monitor.scala 670:37]
  assign _GEN_30 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_29; // @[Monitor.scala 670:37]
  assign _T_1041 = io_in_d_bits_opcode == _GEN_30; // @[Monitor.scala 670:37]
  assign _GEN_37 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_28; // @[Monitor.scala 670:96]
  assign _GEN_38 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_37; // @[Monitor.scala 670:96]
  assign _T_1043 = io_in_d_bits_opcode == _GEN_38; // @[Monitor.scala 670:96]
  assign _T_1044 = _T_1041 | _T_1043; // @[Monitor.scala 670:71]
  assign _T_1047 = _T_781 | _T_781; // @[Monitor.scala 671:99]
  assign _T_1048 = io_in_a_valid & _T_1047; // @[Monitor.scala 671:34]
  assign _T_1049 = _T_1044 | _T_1048; // @[Monitor.scala 671:15]
  assign _T_1051 = _T_1049 | reset; // @[Monitor.scala 51:11]
  assign a_size_lookup = _T_985[7:0]; // @[Monitor.scala 636:19]
  assign _GEN_60 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 673:34]
  assign _T_1053 = _GEN_60 == a_size_lookup; // @[Monitor.scala 673:34]
  assign _T_1056 = _T_1053 | _T_1034; // @[Monitor.scala 673:53]
  assign _T_1058 = _T_1056 | reset; // @[Monitor.scala 51:11]
  assign _T_1061 = _T_1008 & a_first; // @[Monitor.scala 675:36]
  assign _T_1062 = _T_1061 & io_in_a_valid; // @[Monitor.scala 675:47]
  assign _T_1066 = _T_1062 & ~_T_687; // @[Monitor.scala 675:116]
  assign _T_1070 = io_in_a_ready | reset; // @[Monitor.scala 51:11]
  assign a_set = _GEN_15[0]; // @[Monitor.scala 647:13]
  assign d_clr = _GEN_20[0]; // @[Monitor.scala 664:13]
  assign _T_1072 = a_set != d_clr; // @[Monitor.scala 680:20]
  assign _T_1073 = |a_set; // @[Monitor.scala 680:40]
  assign _T_1075 = _T_1072 | ~_T_1073; // @[Monitor.scala 680:30]
  assign _T_1077 = _T_1075 | reset; // @[Monitor.scala 51:11]
  assign _T_1079 = inflight | a_set; // @[Monitor.scala 683:27]
  assign _T_1081 = _T_1079 & ~d_clr; // @[Monitor.scala 683:36]
  assign a_opcodes_set = _GEN_18[3:0]; // @[Monitor.scala 650:21]
  assign _T_1082 = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 684:43]
  assign d_opcodes_clr = _GEN_21[3:0]; // @[Monitor.scala 665:21]
  assign _T_1084 = _T_1082 & ~d_opcodes_clr; // @[Monitor.scala 684:60]
  assign a_sizes_set = _GEN_19[7:0]; // @[Monitor.scala 651:19]
  assign _T_1085 = inflight_sizes | a_sizes_set; // @[Monitor.scala 685:39]
  assign d_sizes_clr = _GEN_22[7:0]; // @[Monitor.scala 666:19]
  assign _T_1087 = _T_1085 & ~d_sizes_clr; // @[Monitor.scala 685:54]
  assign _GEN_61 = io_in_d_valid & _T_687; // @[Monitor.scala 51:11]
  assign _GEN_69 = io_in_d_valid & _T_707; // @[Monitor.scala 51:11]
  assign _GEN_77 = io_in_d_valid & _T_735; // @[Monitor.scala 51:11]
  assign _GEN_85 = io_in_d_valid & _T_764; // @[Monitor.scala 51:11]
  assign _GEN_89 = io_in_d_valid & _T_781; // @[Monitor.scala 51:11]
  assign _GEN_93 = io_in_d_valid & _T_799; // @[Monitor.scala 51:11]
  assign TLMonitor_36_covSum = 30'h0;
  assign io_covSum = TLMonitor_36_covSum;
  assign stopEn0 = io_in_a_valid & ~_T_288;
  assign stopEn1 = io_in_a_valid & ~_T_140;
  assign stopEn2 = io_in_d_valid & ~_T_682;
  assign stopEn3 = _GEN_61 & ~_T_693;
  assign stopEn4 = _GEN_61 & ~_T_697;
  assign stopEn5 = _GEN_61 & ~_T_701;
  assign stopEn6 = _GEN_61 & ~_T_705;
  assign stopEn7 = _GEN_69 & ~_T_693;
  assign stopEn8 = _GEN_69 & ~_T_720;
  assign stopEn9 = _GEN_69 & ~_T_724;
  assign stopEn10 = _GEN_69 & ~_T_701;
  assign stopEn11 = _GEN_77 & ~_T_693;
  assign stopEn12 = _GEN_77 & ~_T_720;
  assign stopEn13 = _GEN_77 & ~_T_724;
  assign stopEn14 = _GEN_77 & ~_T_757;
  assign stopEn15 = _GEN_85 & ~_T_697;
  assign stopEn16 = _GEN_85 & ~_T_701;
  assign stopEn17 = _GEN_89 & ~_T_697;
  assign stopEn18 = _GEN_89 & ~_T_757;
  assign stopEn19 = _GEN_93 & ~_T_697;
  assign stopEn20 = _GEN_93 & ~_T_701;
  assign stopEn21 = _T_857 & ~_T_876;
  assign stopEn22 = _T_906 & ~_T_909;
  assign stopEn23 = _T_906 & ~_T_913;
  assign stopEn24 = _T_906 & ~_T_917;
  assign stopEn25 = _T_906 & ~_T_925;
  assign stopEn26 = _T_906 & ~_T_929;
  assign stopEn27 = _T_989 & ~_T_1004;
  assign stopEn28 = _T_1011 & ~_T_1038;
  assign stopEn29 = _T_1011 & ~_T_1051;
  assign stopEn30 = _T_1011 & ~_T_1058;
  assign stopEn31 = _T_1066 & ~_T_1070;
  assign stopEn32 = ~_T_1077;
  assign TLMonitor_36_or15 = stopEn0 | stopEn1;
  assign TLMonitor_36_or16 = stopEn2 | stopEn3;
  assign TLMonitor_36_or7 = TLMonitor_36_or15 | TLMonitor_36_or16;
  assign TLMonitor_36_or17 = stopEn4 | stopEn5;
  assign TLMonitor_36_or18 = stopEn6 | stopEn7;
  assign TLMonitor_36_or8 = TLMonitor_36_or17 | TLMonitor_36_or18;
  assign TLMonitor_36_or3 = TLMonitor_36_or7 | TLMonitor_36_or8;
  assign TLMonitor_36_or19 = stopEn8 | stopEn9;
  assign TLMonitor_36_or20 = stopEn10 | stopEn11;
  assign TLMonitor_36_or9 = TLMonitor_36_or19 | TLMonitor_36_or20;
  assign TLMonitor_36_or21 = stopEn12 | stopEn13;
  assign TLMonitor_36_or22 = stopEn14 | stopEn15;
  assign TLMonitor_36_or10 = TLMonitor_36_or21 | TLMonitor_36_or22;
  assign TLMonitor_36_or4 = TLMonitor_36_or9 | TLMonitor_36_or10;
  assign TLMonitor_36_or1 = TLMonitor_36_or3 | TLMonitor_36_or4;
  assign TLMonitor_36_or23 = stopEn16 | stopEn17;
  assign TLMonitor_36_or24 = stopEn18 | stopEn19;
  assign TLMonitor_36_or11 = TLMonitor_36_or23 | TLMonitor_36_or24;
  assign TLMonitor_36_or25 = stopEn20 | stopEn21;
  assign TLMonitor_36_or26 = stopEn22 | stopEn23;
  assign TLMonitor_36_or12 = TLMonitor_36_or25 | TLMonitor_36_or26;
  assign TLMonitor_36_or5 = TLMonitor_36_or11 | TLMonitor_36_or12;
  assign TLMonitor_36_or27 = stopEn24 | stopEn25;
  assign TLMonitor_36_or28 = stopEn26 | stopEn27;
  assign TLMonitor_36_or13 = TLMonitor_36_or27 | TLMonitor_36_or28;
  assign TLMonitor_36_or29 = stopEn28 | stopEn29;
  assign TLMonitor_36_or62 = stopEn31 | stopEn32;
  assign TLMonitor_36_or30 = stopEn30 | TLMonitor_36_or62;
  assign TLMonitor_36_or14 = TLMonitor_36_or29 | TLMonitor_36_or30;
  assign TLMonitor_36_or6 = TLMonitor_36_or13 | TLMonitor_36_or14;
  assign TLMonitor_36_or2 = TLMonitor_36_or5 | TLMonitor_36_or6;
  assign TLMonitor_36_or0 = TLMonitor_36_or1 | TLMonitor_36_or2;
  assign metaAssert = TLMonitor_36_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_840 = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_855 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_888 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_899 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_900 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_901 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_903 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_904 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  inflight = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  inflight_opcodes = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  inflight_sizes = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_942 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_960 = _RAND_12[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  TLMonitor_36_metaAssert = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_840 <= 9'h0;
    end else if (reset) begin
      _T_840 <= 9'h0;
    end else if (_T_831) begin
      if (_T_843) begin
        _T_840 <= 9'h0;
      end else begin
        _T_840 <= _T_842;
      end
    end
    if (metaReset) begin
      _T_855 <= 32'h0;
    end else if (_T_879) begin
      _T_855 <= io_in_a_bits_address;
    end
    if (metaReset) begin
      _T_888 <= 9'h0;
    end else if (reset) begin
      _T_888 <= 9'h0;
    end else if (io_in_d_valid) begin
      if (_T_891) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_888 <= _T_885;
        end else begin
          _T_888 <= 9'h0;
        end
      end else begin
        _T_888 <= _T_890;
      end
    end
    if (metaReset) begin
      _T_899 <= 3'h0;
    end else if (_T_932) begin
      _T_899 <= io_in_d_bits_opcode;
    end
    if (metaReset) begin
      _T_900 <= 2'h0;
    end else if (_T_932) begin
      _T_900 <= io_in_d_bits_param;
    end
    if (metaReset) begin
      _T_901 <= 4'h0;
    end else if (_T_932) begin
      _T_901 <= io_in_d_bits_size;
    end
    if (metaReset) begin
      _T_903 <= 2'h0;
    end else if (_T_932) begin
      _T_903 <= io_in_d_bits_sink;
    end
    if (metaReset) begin
      _T_904 <= 1'h0;
    end else if (_T_932) begin
      _T_904 <= io_in_d_bits_denied;
    end
    if (metaReset) begin
      inflight <= 1'h0;
    end else if (reset) begin
      inflight <= 1'h0;
    end else begin
      inflight <= _T_1081;
    end
    if (metaReset) begin
      inflight_opcodes <= 4'h0;
    end else if (reset) begin
      inflight_opcodes <= 4'h0;
    end else begin
      inflight_opcodes <= _T_1084;
    end
    if (metaReset) begin
      inflight_sizes <= 8'h0;
    end else if (reset) begin
      inflight_sizes <= 8'h0;
    end else begin
      inflight_sizes <= _T_1087;
    end
    if (metaReset) begin
      _T_942 <= 9'h0;
    end else if (reset) begin
      _T_942 <= 9'h0;
    end else if (_T_831) begin
      if (a_first) begin
        _T_942 <= 9'h0;
      end else begin
        _T_942 <= _T_944;
      end
    end
    if (metaReset) begin
      _T_960 <= 9'h0;
    end else if (reset) begin
      _T_960 <= 9'h0;
    end else if (io_in_d_valid) begin
      if (d_first) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_960 <= _T_885;
        end else begin
          _T_960 <= 9'h0;
        end
      end else begin
        _T_960 <= _T_962;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & ~_T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type which is unexpected using diplomatic parameters\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at Frontend.scala:353:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & ~_T_288) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & ~_T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at Frontend.scala:353:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & ~_T_140) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~_T_682) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~_T_682) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_61 & ~_T_693) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_61 & ~_T_693) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_61 & ~_T_697) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_61 & ~_T_697) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_61 & ~_T_701) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_61 & ~_T_701) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_61 & ~_T_705) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_61 & ~_T_705) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & ~_T_693) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & ~_T_693) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & ~_T_720) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & ~_T_720) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & ~_T_724) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & ~_T_724) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & ~_T_701) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & ~_T_701) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_77 & ~_T_693) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_77 & ~_T_693) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_77 & ~_T_720) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_77 & ~_T_720) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_77 & ~_T_724) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_77 & ~_T_724) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_77 & ~_T_757) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_77 & ~_T_757) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & ~_T_697) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & ~_T_697) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & ~_T_701) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & ~_T_701) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_89 & ~_T_697) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_89 & ~_T_697) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_89 & ~_T_757) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_89 & ~_T_757) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & ~_T_697) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & ~_T_697) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & ~_T_701) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & ~_T_701) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_857 & ~_T_876) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at Frontend.scala:353:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_857 & ~_T_876) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_906 & ~_T_909) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_906 & ~_T_909) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_906 & ~_T_913) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_906 & ~_T_913) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_906 & ~_T_917) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_906 & ~_T_917) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_906 & ~_T_925) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_906 & ~_T_925) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_906 & ~_T_929) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_906 & ~_T_929) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_989 & ~_T_1004) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at Frontend.scala:353:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_989 & ~_T_1004) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1011 & ~_T_1038) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1011 & ~_T_1038) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1011 & ~_T_1051) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1011 & ~_T_1051) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1011 & ~_T_1058) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1011 & ~_T_1058) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1066 & ~_T_1070) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1066 & ~_T_1070) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1077) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at Frontend.scala:353:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1077) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    if (metaReset) begin
      TLMonitor_36_metaAssert <= 1'h0;
    end else begin
      TLMonitor_36_metaAssert <= TLMonitor_36_metaAssert | TLMonitor_36_or0;
    end
  end
endmodule
module TLB(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [39:0] io_req_bits_vaddr,
  input         io_req_bits_passthrough,
  input  [1:0]  io_req_bits_size,
  input  [4:0]  io_req_bits_cmd,
  output        io_resp_miss,
  output [31:0] io_resp_paddr,
  output        io_resp_pf_ld,
  output        io_resp_pf_st,
  output        io_resp_ae_ld,
  output        io_resp_ae_st,
  output        io_resp_ma_ld,
  output        io_resp_ma_st,
  output        io_resp_cacheable,
  input         io_sfence_valid,
  input         io_sfence_bits_rs1,
  input         io_sfence_bits_rs2,
  input  [38:0] io_sfence_bits_addr,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input         io_ptw_status_debug,
  input  [1:0]  io_ptw_status_dprv,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [19:0] OptimizationBarrier_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_metaAssert; // @[package.scala 236:25]
  wire [1:0] pmp_io_prv; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_0_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_0_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_1_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_1_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_2_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_2_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_3_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_3_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_4_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_4_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_5_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_5_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_6_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_6_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_7_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_7_mask; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_addr; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_size; // @[TLB.scala 190:19]
  wire  pmp_io_r; // @[TLB.scala 190:19]
  wire  pmp_io_w; // @[TLB.scala 190:19]
  wire  pmp_io_x; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_covSum; // @[TLB.scala 190:19]
  wire  pmp_metaAssert; // @[TLB.scala 190:19]
  wire [19:0] OptimizationBarrier_1_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_1_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_1_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_2_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_2_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_2_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_3_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_3_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_3_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_4_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_4_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_4_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_5_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_5_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_5_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_6_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_6_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_6_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_7_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_7_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_7_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_8_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_8_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_8_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_9_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_9_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_9_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_10_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_10_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_10_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_11_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_11_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_11_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_12_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_12_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_12_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_13_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_13_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_13_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_14_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_14_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_14_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_15_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_15_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_15_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_16_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_16_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_16_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_17_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_17_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_17_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_18_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_18_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_18_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_19_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_19_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_19_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_20_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_20_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_20_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_21_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_21_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_21_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_22_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_22_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_22_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_23_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_23_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_23_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_24_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_24_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_24_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_25_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_25_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_25_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_26_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_26_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_26_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_27_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_27_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_27_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_28_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_28_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_28_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_29_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_29_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_29_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_30_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_30_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_30_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_31_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_31_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_31_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_32_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_32_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_32_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_33_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_33_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_33_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_34_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_34_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_34_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_35_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_35_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_35_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_36_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_36_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_36_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_37_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_37_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_37_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_38_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_38_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_38_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_metaAssert; // @[package.scala 236:25]
  reg [26:0] sectored_entries_0_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_0;
  reg [34:0] sectored_entries_0_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_1;
  reg [34:0] sectored_entries_0_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_2;
  reg [34:0] sectored_entries_0_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_3;
  reg [34:0] sectored_entries_0_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_4;
  reg  sectored_entries_0_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_5;
  reg  sectored_entries_0_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_6;
  reg  sectored_entries_0_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_7;
  reg  sectored_entries_0_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_8;
  reg [26:0] sectored_entries_1_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_9;
  reg [34:0] sectored_entries_1_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_10;
  reg [34:0] sectored_entries_1_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_11;
  reg [34:0] sectored_entries_1_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_12;
  reg [34:0] sectored_entries_1_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_13;
  reg  sectored_entries_1_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_14;
  reg  sectored_entries_1_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_15;
  reg  sectored_entries_1_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_16;
  reg  sectored_entries_1_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_17;
  reg [26:0] sectored_entries_2_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_18;
  reg [34:0] sectored_entries_2_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_19;
  reg [34:0] sectored_entries_2_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_20;
  reg [34:0] sectored_entries_2_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_21;
  reg [34:0] sectored_entries_2_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_22;
  reg  sectored_entries_2_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_23;
  reg  sectored_entries_2_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_24;
  reg  sectored_entries_2_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_25;
  reg  sectored_entries_2_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_26;
  reg [26:0] sectored_entries_3_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_27;
  reg [34:0] sectored_entries_3_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_28;
  reg [34:0] sectored_entries_3_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_29;
  reg [34:0] sectored_entries_3_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_30;
  reg [34:0] sectored_entries_3_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_31;
  reg  sectored_entries_3_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_32;
  reg  sectored_entries_3_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_33;
  reg  sectored_entries_3_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_34;
  reg  sectored_entries_3_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_35;
  reg [26:0] sectored_entries_4_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_36;
  reg [34:0] sectored_entries_4_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_37;
  reg [34:0] sectored_entries_4_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_38;
  reg [34:0] sectored_entries_4_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_39;
  reg [34:0] sectored_entries_4_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_40;
  reg  sectored_entries_4_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_41;
  reg  sectored_entries_4_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_42;
  reg  sectored_entries_4_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_43;
  reg  sectored_entries_4_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_44;
  reg [26:0] sectored_entries_5_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_45;
  reg [34:0] sectored_entries_5_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_46;
  reg [34:0] sectored_entries_5_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_47;
  reg [34:0] sectored_entries_5_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_48;
  reg [34:0] sectored_entries_5_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_49;
  reg  sectored_entries_5_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_50;
  reg  sectored_entries_5_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_51;
  reg  sectored_entries_5_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_52;
  reg  sectored_entries_5_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_53;
  reg [26:0] sectored_entries_6_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_54;
  reg [34:0] sectored_entries_6_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_55;
  reg [34:0] sectored_entries_6_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_56;
  reg [34:0] sectored_entries_6_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_57;
  reg [34:0] sectored_entries_6_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_58;
  reg  sectored_entries_6_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_59;
  reg  sectored_entries_6_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_60;
  reg  sectored_entries_6_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_61;
  reg  sectored_entries_6_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_62;
  reg [26:0] sectored_entries_7_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_63;
  reg [34:0] sectored_entries_7_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_64;
  reg [34:0] sectored_entries_7_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_65;
  reg [34:0] sectored_entries_7_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_66;
  reg [34:0] sectored_entries_7_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_67;
  reg  sectored_entries_7_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_68;
  reg  sectored_entries_7_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_69;
  reg  sectored_entries_7_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_70;
  reg  sectored_entries_7_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_71;
  reg [1:0] superpage_entries_0_level; // @[TLB.scala 163:30]
  reg [31:0] _RAND_72;
  reg [26:0] superpage_entries_0_tag; // @[TLB.scala 163:30]
  reg [31:0] _RAND_73;
  reg [34:0] superpage_entries_0_data_0; // @[TLB.scala 163:30]
  reg [63:0] _RAND_74;
  reg  superpage_entries_0_valid_0; // @[TLB.scala 163:30]
  reg [31:0] _RAND_75;
  reg [1:0] superpage_entries_1_level; // @[TLB.scala 163:30]
  reg [31:0] _RAND_76;
  reg [26:0] superpage_entries_1_tag; // @[TLB.scala 163:30]
  reg [31:0] _RAND_77;
  reg [34:0] superpage_entries_1_data_0; // @[TLB.scala 163:30]
  reg [63:0] _RAND_78;
  reg  superpage_entries_1_valid_0; // @[TLB.scala 163:30]
  reg [31:0] _RAND_79;
  reg [1:0] superpage_entries_2_level; // @[TLB.scala 163:30]
  reg [31:0] _RAND_80;
  reg [26:0] superpage_entries_2_tag; // @[TLB.scala 163:30]
  reg [31:0] _RAND_81;
  reg [34:0] superpage_entries_2_data_0; // @[TLB.scala 163:30]
  reg [63:0] _RAND_82;
  reg  superpage_entries_2_valid_0; // @[TLB.scala 163:30]
  reg [31:0] _RAND_83;
  reg [1:0] superpage_entries_3_level; // @[TLB.scala 163:30]
  reg [31:0] _RAND_84;
  reg [26:0] superpage_entries_3_tag; // @[TLB.scala 163:30]
  reg [31:0] _RAND_85;
  reg [34:0] superpage_entries_3_data_0; // @[TLB.scala 163:30]
  reg [63:0] _RAND_86;
  reg  superpage_entries_3_valid_0; // @[TLB.scala 163:30]
  reg [31:0] _RAND_87;
  reg [1:0] special_entry_level; // @[TLB.scala 164:56]
  reg [31:0] _RAND_88;
  reg [26:0] special_entry_tag; // @[TLB.scala 164:56]
  reg [31:0] _RAND_89;
  reg [34:0] special_entry_data_0; // @[TLB.scala 164:56]
  reg [63:0] _RAND_90;
  reg  special_entry_valid_0; // @[TLB.scala 164:56]
  reg [31:0] _RAND_91;
  reg [1:0] state; // @[TLB.scala 169:18]
  reg [31:0] _RAND_92;
  reg [26:0] r_refill_tag; // @[TLB.scala 170:25]
  reg [31:0] _RAND_93;
  reg [1:0] r_superpage_repl_addr; // @[TLB.scala 171:34]
  reg [31:0] _RAND_94;
  reg [2:0] r_sectored_repl_addr; // @[TLB.scala 172:33]
  reg [31:0] _RAND_95;
  reg [2:0] r_sectored_hit_addr; // @[TLB.scala 173:32]
  reg [31:0] _RAND_96;
  reg  r_sectored_hit; // @[TLB.scala 174:27]
  reg [31:0] _RAND_97;
  wire  priv_s; // @[TLB.scala 177:20]
  wire  priv_uses_vm; // @[TLB.scala 178:27]
  wire  _T_2; // @[TLB.scala 179:83]
  wire  vm_enabled; // @[TLB.scala 179:99]
  wire [26:0] vpn; // @[TLB.scala 182:30]
  wire [19:0] refill_ppn; // @[TLB.scala 183:44]
  wire  _T_4; // @[package.scala 15:47]
  wire  _T_5; // @[package.scala 15:47]
  wire  _T_6; // @[package.scala 64:59]
  wire  invalidate_refill; // @[TLB.scala 185:88]
  wire  _T_27; // @[TLB.scala 108:28]
  wire [26:0] _T_29; // @[TLB.scala 109:28]
  wire [26:0] _GEN_983; // @[TLB.scala 109:47]
  wire [26:0] _T_30; // @[TLB.scala 109:47]
  wire  _T_33; // @[TLB.scala 108:28]
  wire [26:0] _T_35; // @[TLB.scala 109:28]
  wire [26:0] _T_36; // @[TLB.scala 109:47]
  wire [19:0] _T_38; // @[Cat.scala 29:58]
  wire [27:0] _T_40; // @[TLB.scala 187:20]
  wire [27:0] mpu_ppn; // @[TLB.scala 186:20]
  wire [39:0] mpu_physaddr; // @[Cat.scala 29:58]
  wire  _T_42; // @[TLB.scala 189:56]
  wire [2:0] _T_44; // @[Cat.scala 29:58]
  wire [2:0] mpu_priv; // @[TLB.scala 189:27]
  wire [39:0] _T_45; // @[Parameters.scala 137:31]
  wire [40:0] _T_46; // @[Parameters.scala 137:49]
  wire [40:0] _T_48; // @[Parameters.scala 137:52]
  wire  _T_49; // @[Parameters.scala 137:67]
  wire [39:0] _T_50; // @[Parameters.scala 137:31]
  wire [40:0] _T_51; // @[Parameters.scala 137:49]
  wire [40:0] _T_53; // @[Parameters.scala 137:52]
  wire  _T_54; // @[Parameters.scala 137:67]
  wire [39:0] _T_55; // @[Parameters.scala 137:31]
  wire [40:0] _T_56; // @[Parameters.scala 137:49]
  wire [40:0] _T_58; // @[Parameters.scala 137:52]
  wire  _T_59; // @[Parameters.scala 137:67]
  wire [40:0] _T_61; // @[Parameters.scala 137:49]
  wire [40:0] _T_63; // @[Parameters.scala 137:52]
  wire  _T_64; // @[Parameters.scala 137:67]
  wire [39:0] _T_65; // @[Parameters.scala 137:31]
  wire [40:0] _T_66; // @[Parameters.scala 137:49]
  wire [40:0] _T_68; // @[Parameters.scala 137:52]
  wire  _T_69; // @[Parameters.scala 137:67]
  wire [39:0] _T_70; // @[Parameters.scala 137:31]
  wire [40:0] _T_71; // @[Parameters.scala 137:49]
  wire [40:0] _T_73; // @[Parameters.scala 137:52]
  wire  _T_74; // @[Parameters.scala 137:67]
  wire [39:0] _T_75; // @[Parameters.scala 137:31]
  wire [40:0] _T_76; // @[Parameters.scala 137:49]
  wire [40:0] _T_78; // @[Parameters.scala 137:52]
  wire  _T_79; // @[Parameters.scala 137:67]
  wire  _T_81; // @[TLB.scala 195:67]
  wire  _T_82; // @[TLB.scala 195:67]
  wire  _T_83; // @[TLB.scala 195:67]
  wire  _T_84; // @[TLB.scala 195:67]
  wire  _T_85; // @[TLB.scala 195:67]
  wire  legal_address; // @[TLB.scala 195:67]
  wire [40:0] _T_94; // @[Parameters.scala 137:52]
  wire  _T_95; // @[Parameters.scala 137:67]
  wire  cacheable; // @[TLB.scala 197:19]
  wire [39:0] _T_155; // @[Parameters.scala 137:31]
  wire [40:0] _T_156; // @[Parameters.scala 137:49]
  wire [40:0] _T_158; // @[Parameters.scala 137:52]
  wire  _T_159; // @[Parameters.scala 137:67]
  wire [40:0] _T_172; // @[Parameters.scala 137:52]
  wire  _T_173; // @[Parameters.scala 137:67]
  wire  _T_180; // @[TLBPermissions.scala 82:66]
  wire  _T_193; // @[TLB.scala 200:39]
  wire  deny_access_to_debug; // @[TLB.scala 200:48]
  wire  _T_206; // @[TLB.scala 201:41]
  wire  prot_r; // @[TLB.scala 201:66]
  wire [39:0] _T_217; // @[Parameters.scala 137:31]
  wire [40:0] _T_218; // @[Parameters.scala 137:49]
  wire [40:0] _T_220; // @[Parameters.scala 137:52]
  wire  _T_221; // @[Parameters.scala 137:67]
  wire [40:0] _T_225; // @[Parameters.scala 137:52]
  wire  _T_226; // @[Parameters.scala 137:67]
  wire  _T_228; // @[Parameters.scala 549:89]
  wire  _T_229; // @[Parameters.scala 549:89]
  wire  _T_239; // @[TLB.scala 197:19]
  wire  _T_241; // @[TLB.scala 202:45]
  wire  prot_w; // @[TLB.scala 202:70]
  wire  prot_al; // @[TLB.scala 197:19]
  wire [40:0] _T_341; // @[Parameters.scala 137:52]
  wire  _T_342; // @[Parameters.scala 137:67]
  wire  _T_353; // @[Parameters.scala 549:89]
  wire  _T_354; // @[Parameters.scala 549:89]
  wire  _T_370; // @[TLB.scala 197:19]
  wire  _T_372; // @[TLB.scala 206:40]
  wire  prot_x; // @[TLB.scala 206:65]
  wire [40:0] _T_393; // @[Parameters.scala 137:52]
  wire  _T_394; // @[Parameters.scala 137:67]
  wire [40:0] _T_398; // @[Parameters.scala 137:52]
  wire  _T_399; // @[Parameters.scala 137:67]
  wire  _T_410; // @[Parameters.scala 549:89]
  wire  _T_411; // @[Parameters.scala 549:89]
  wire  _T_412; // @[Parameters.scala 549:89]
  wire  prot_eff; // @[TLB.scala 197:19]
  wire  _T_417; // @[package.scala 64:59]
  wire  _T_418; // @[package.scala 64:59]
  wire  _T_419; // @[package.scala 64:59]
  wire [26:0] _T_420; // @[TLB.scala 88:41]
  wire  _T_422; // @[TLB.scala 88:66]
  wire  sector_hits_0; // @[TLB.scala 87:40]
  wire  _T_423; // @[package.scala 64:59]
  wire  _T_424; // @[package.scala 64:59]
  wire  _T_425; // @[package.scala 64:59]
  wire [26:0] _T_426; // @[TLB.scala 88:41]
  wire  _T_428; // @[TLB.scala 88:66]
  wire  sector_hits_1; // @[TLB.scala 87:40]
  wire  _T_429; // @[package.scala 64:59]
  wire  _T_430; // @[package.scala 64:59]
  wire  _T_431; // @[package.scala 64:59]
  wire [26:0] _T_432; // @[TLB.scala 88:41]
  wire  _T_434; // @[TLB.scala 88:66]
  wire  sector_hits_2; // @[TLB.scala 87:40]
  wire  _T_435; // @[package.scala 64:59]
  wire  _T_436; // @[package.scala 64:59]
  wire  _T_437; // @[package.scala 64:59]
  wire [26:0] _T_438; // @[TLB.scala 88:41]
  wire  _T_440; // @[TLB.scala 88:66]
  wire  sector_hits_3; // @[TLB.scala 87:40]
  wire  _T_441; // @[package.scala 64:59]
  wire  _T_442; // @[package.scala 64:59]
  wire  _T_443; // @[package.scala 64:59]
  wire [26:0] _T_444; // @[TLB.scala 88:41]
  wire  _T_446; // @[TLB.scala 88:66]
  wire  sector_hits_4; // @[TLB.scala 87:40]
  wire  _T_447; // @[package.scala 64:59]
  wire  _T_448; // @[package.scala 64:59]
  wire  _T_449; // @[package.scala 64:59]
  wire [26:0] _T_450; // @[TLB.scala 88:41]
  wire  _T_452; // @[TLB.scala 88:66]
  wire  sector_hits_5; // @[TLB.scala 87:40]
  wire  _T_453; // @[package.scala 64:59]
  wire  _T_454; // @[package.scala 64:59]
  wire  _T_455; // @[package.scala 64:59]
  wire [26:0] _T_456; // @[TLB.scala 88:41]
  wire  _T_458; // @[TLB.scala 88:66]
  wire  sector_hits_6; // @[TLB.scala 87:40]
  wire  _T_459; // @[package.scala 64:59]
  wire  _T_460; // @[package.scala 64:59]
  wire  _T_461; // @[package.scala 64:59]
  wire [26:0] _T_462; // @[TLB.scala 88:41]
  wire  _T_464; // @[TLB.scala 88:66]
  wire  sector_hits_7; // @[TLB.scala 87:40]
  wire  _T_469; // @[TLB.scala 95:77]
  wire  _T_471; // @[TLB.scala 95:29]
  wire  _T_472; // @[TLB.scala 94:28]
  wire  _T_476; // @[TLB.scala 95:77]
  wire  _T_477; // @[TLB.scala 95:40]
  wire  superpage_hits_0; // @[TLB.scala 95:29]
  wire  _T_489; // @[TLB.scala 95:77]
  wire  _T_491; // @[TLB.scala 95:29]
  wire  _T_492; // @[TLB.scala 94:28]
  wire  _T_496; // @[TLB.scala 95:77]
  wire  _T_497; // @[TLB.scala 95:40]
  wire  superpage_hits_1; // @[TLB.scala 95:29]
  wire  _T_509; // @[TLB.scala 95:77]
  wire  _T_511; // @[TLB.scala 95:29]
  wire  _T_512; // @[TLB.scala 94:28]
  wire  _T_516; // @[TLB.scala 95:77]
  wire  _T_517; // @[TLB.scala 95:40]
  wire  superpage_hits_2; // @[TLB.scala 95:29]
  wire  _T_529; // @[TLB.scala 95:77]
  wire  _T_531; // @[TLB.scala 95:29]
  wire  _T_532; // @[TLB.scala 94:28]
  wire  _T_536; // @[TLB.scala 95:77]
  wire  _T_537; // @[TLB.scala 95:40]
  wire  superpage_hits_3; // @[TLB.scala 95:29]
  wire  _GEN_1; // @[TLB.scala 100:18]
  wire  _GEN_2; // @[TLB.scala 100:18]
  wire  _GEN_3; // @[TLB.scala 100:18]
  wire  _T_549; // @[TLB.scala 100:18]
  wire  hitsVec_0; // @[TLB.scala 211:44]
  wire  _GEN_5; // @[TLB.scala 100:18]
  wire  _GEN_6; // @[TLB.scala 100:18]
  wire  _GEN_7; // @[TLB.scala 100:18]
  wire  _T_554; // @[TLB.scala 100:18]
  wire  hitsVec_1; // @[TLB.scala 211:44]
  wire  _GEN_9; // @[TLB.scala 100:18]
  wire  _GEN_10; // @[TLB.scala 100:18]
  wire  _GEN_11; // @[TLB.scala 100:18]
  wire  _T_559; // @[TLB.scala 100:18]
  wire  hitsVec_2; // @[TLB.scala 211:44]
  wire  _GEN_13; // @[TLB.scala 100:18]
  wire  _GEN_14; // @[TLB.scala 100:18]
  wire  _GEN_15; // @[TLB.scala 100:18]
  wire  _T_564; // @[TLB.scala 100:18]
  wire  hitsVec_3; // @[TLB.scala 211:44]
  wire  _GEN_17; // @[TLB.scala 100:18]
  wire  _GEN_18; // @[TLB.scala 100:18]
  wire  _GEN_19; // @[TLB.scala 100:18]
  wire  _T_569; // @[TLB.scala 100:18]
  wire  hitsVec_4; // @[TLB.scala 211:44]
  wire  _GEN_21; // @[TLB.scala 100:18]
  wire  _GEN_22; // @[TLB.scala 100:18]
  wire  _GEN_23; // @[TLB.scala 100:18]
  wire  _T_574; // @[TLB.scala 100:18]
  wire  hitsVec_5; // @[TLB.scala 211:44]
  wire  _GEN_25; // @[TLB.scala 100:18]
  wire  _GEN_26; // @[TLB.scala 100:18]
  wire  _GEN_27; // @[TLB.scala 100:18]
  wire  _T_579; // @[TLB.scala 100:18]
  wire  hitsVec_6; // @[TLB.scala 211:44]
  wire  _GEN_29; // @[TLB.scala 100:18]
  wire  _GEN_30; // @[TLB.scala 100:18]
  wire  _GEN_31; // @[TLB.scala 100:18]
  wire  _T_584; // @[TLB.scala 100:18]
  wire  hitsVec_7; // @[TLB.scala 211:44]
  wire  hitsVec_8; // @[TLB.scala 211:44]
  wire  hitsVec_9; // @[TLB.scala 211:44]
  wire  hitsVec_10; // @[TLB.scala 211:44]
  wire  hitsVec_11; // @[TLB.scala 211:44]
  wire  _T_673; // @[TLB.scala 95:77]
  wire  _T_675; // @[TLB.scala 95:29]
  wire  _T_680; // @[TLB.scala 95:77]
  wire  _T_681; // @[TLB.scala 95:40]
  wire  _T_682; // @[TLB.scala 95:29]
  wire  _T_687; // @[TLB.scala 95:77]
  wire  _T_688; // @[TLB.scala 95:40]
  wire  _T_689; // @[TLB.scala 95:29]
  wire  hitsVec_12; // @[TLB.scala 211:44]
  wire [5:0] _T_694; // @[Cat.scala 29:58]
  wire [12:0] real_hits; // @[Cat.scala 29:58]
  wire [13:0] hits; // @[Cat.scala 29:58]
  wire [34:0] _GEN_33;
  wire [34:0] _GEN_34;
  wire [34:0] _GEN_35;
  wire [34:0] _GEN_37;
  wire [34:0] _GEN_38;
  wire [34:0] _GEN_39;
  wire [34:0] _GEN_41;
  wire [34:0] _GEN_42;
  wire [34:0] _GEN_43;
  wire [34:0] _GEN_45;
  wire [34:0] _GEN_46;
  wire [34:0] _GEN_47;
  wire [34:0] _GEN_49;
  wire [34:0] _GEN_50;
  wire [34:0] _GEN_51;
  wire [34:0] _GEN_53;
  wire [34:0] _GEN_54;
  wire [34:0] _GEN_55;
  wire [34:0] _GEN_57;
  wire [34:0] _GEN_58;
  wire [34:0] _GEN_59;
  wire [34:0] _GEN_61;
  wire [34:0] _GEN_62;
  wire [34:0] _GEN_63;
  wire [26:0] _T_876; // @[TLB.scala 109:28]
  wire [26:0] _GEN_985; // @[TLB.scala 109:47]
  wire [26:0] _T_877; // @[TLB.scala 109:47]
  wire [26:0] _T_883; // @[TLB.scala 109:47]
  wire [19:0] _T_885; // @[Cat.scala 29:58]
  wire [26:0] _T_907; // @[TLB.scala 109:28]
  wire [26:0] _GEN_987; // @[TLB.scala 109:47]
  wire [26:0] _T_908; // @[TLB.scala 109:47]
  wire [26:0] _T_914; // @[TLB.scala 109:47]
  wire [19:0] _T_916; // @[Cat.scala 29:58]
  wire [26:0] _T_938; // @[TLB.scala 109:28]
  wire [26:0] _GEN_989; // @[TLB.scala 109:47]
  wire [26:0] _T_939; // @[TLB.scala 109:47]
  wire [26:0] _T_945; // @[TLB.scala 109:47]
  wire [19:0] _T_947; // @[Cat.scala 29:58]
  wire [26:0] _T_969; // @[TLB.scala 109:28]
  wire [26:0] _GEN_991; // @[TLB.scala 109:47]
  wire [26:0] _T_970; // @[TLB.scala 109:47]
  wire [26:0] _T_976; // @[TLB.scala 109:47]
  wire [19:0] _T_978; // @[Cat.scala 29:58]
  wire [26:0] _GEN_993; // @[TLB.scala 109:47]
  wire [26:0] _T_1001; // @[TLB.scala 109:47]
  wire [26:0] _T_1007; // @[TLB.scala 109:47]
  wire [19:0] _T_1009; // @[Cat.scala 29:58]
  wire [19:0] _T_1011; // @[Mux.scala 27:72]
  wire [19:0] _T_1012; // @[Mux.scala 27:72]
  wire [19:0] _T_1013; // @[Mux.scala 27:72]
  wire [19:0] _T_1014; // @[Mux.scala 27:72]
  wire [19:0] _T_1015; // @[Mux.scala 27:72]
  wire [19:0] _T_1016; // @[Mux.scala 27:72]
  wire [19:0] _T_1017; // @[Mux.scala 27:72]
  wire [19:0] _T_1018; // @[Mux.scala 27:72]
  wire [19:0] _T_1019; // @[Mux.scala 27:72]
  wire [19:0] _T_1020; // @[Mux.scala 27:72]
  wire [19:0] _T_1021; // @[Mux.scala 27:72]
  wire [19:0] _T_1022; // @[Mux.scala 27:72]
  wire [19:0] _T_1023; // @[Mux.scala 27:72]
  wire [19:0] _T_1024; // @[Mux.scala 27:72]
  wire [19:0] _T_1025; // @[Mux.scala 27:72]
  wire [19:0] _T_1026; // @[Mux.scala 27:72]
  wire [19:0] _T_1027; // @[Mux.scala 27:72]
  wire [19:0] _T_1028; // @[Mux.scala 27:72]
  wire [19:0] _T_1029; // @[Mux.scala 27:72]
  wire [19:0] _T_1030; // @[Mux.scala 27:72]
  wire [19:0] _T_1031; // @[Mux.scala 27:72]
  wire [19:0] _T_1032; // @[Mux.scala 27:72]
  wire [19:0] _T_1033; // @[Mux.scala 27:72]
  wire [19:0] _T_1034; // @[Mux.scala 27:72]
  wire [19:0] _T_1035; // @[Mux.scala 27:72]
  wire [19:0] _T_1036; // @[Mux.scala 27:72]
  wire [19:0] ppn; // @[Mux.scala 27:72]
  wire  _T_1039; // @[TLB.scala 223:25]
  wire  _T_1041; // @[PTW.scala 69:44]
  wire  _T_1042; // @[PTW.scala 69:38]
  wire  _T_1043; // @[PTW.scala 69:32]
  wire  _T_1044; // @[PTW.scala 69:52]
  wire  _T_1045; // @[PTW.scala 73:35]
  wire  _T_1051; // @[PTW.scala 74:35]
  wire  _T_1052; // @[PTW.scala 74:40]
  wire  _T_1058; // @[PTW.scala 75:35]
  wire [7:0] _T_1068; // @[TLB.scala 123:24]
  wire [34:0] _T_1076; // @[TLB.scala 123:24]
  wire  _GEN_64; // @[TLB.scala 240:34]
  wire  _T_1077; // @[TLB.scala 242:40]
  wire  _T_1078; // @[TLB.scala 243:82]
  wire  _GEN_67; // @[TLB.scala 243:89]
  wire  _T_1095; // @[TLB.scala 243:82]
  wire  _GEN_71; // @[TLB.scala 243:89]
  wire  _T_1112; // @[TLB.scala 243:82]
  wire  _GEN_75; // @[TLB.scala 243:89]
  wire  _T_1129; // @[TLB.scala 243:82]
  wire  _GEN_79; // @[TLB.scala 243:89]
  wire [2:0] _T_1146; // @[TLB.scala 248:22]
  wire  _T_1147; // @[TLB.scala 249:65]
  wire  _GEN_81; // @[TLB.scala 250:32]
  wire  _GEN_82; // @[TLB.scala 250:32]
  wire  _GEN_83; // @[TLB.scala 250:32]
  wire  _GEN_84; // @[TLB.scala 250:32]
  wire  _GEN_995; // @[TLB.scala 122:16]
  wire  _GEN_85; // @[TLB.scala 122:16]
  wire  _GEN_996; // @[TLB.scala 122:16]
  wire  _GEN_86; // @[TLB.scala 122:16]
  wire  _GEN_997; // @[TLB.scala 122:16]
  wire  _GEN_87; // @[TLB.scala 122:16]
  wire  _GEN_998; // @[TLB.scala 122:16]
  wire  _GEN_88; // @[TLB.scala 122:16]
  wire  _GEN_93; // @[TLB.scala 252:34]
  wire  _GEN_94; // @[TLB.scala 252:34]
  wire  _GEN_95; // @[TLB.scala 252:34]
  wire  _GEN_96; // @[TLB.scala 252:34]
  wire  _GEN_97; // @[TLB.scala 249:72]
  wire  _GEN_98; // @[TLB.scala 249:72]
  wire  _GEN_99; // @[TLB.scala 249:72]
  wire  _GEN_100; // @[TLB.scala 249:72]
  wire  _T_1165; // @[TLB.scala 249:65]
  wire  _GEN_107; // @[TLB.scala 250:32]
  wire  _GEN_108; // @[TLB.scala 250:32]
  wire  _GEN_109; // @[TLB.scala 250:32]
  wire  _GEN_110; // @[TLB.scala 250:32]
  wire  _GEN_111; // @[TLB.scala 122:16]
  wire  _GEN_112; // @[TLB.scala 122:16]
  wire  _GEN_113; // @[TLB.scala 122:16]
  wire  _GEN_114; // @[TLB.scala 122:16]
  wire  _GEN_119; // @[TLB.scala 252:34]
  wire  _GEN_120; // @[TLB.scala 252:34]
  wire  _GEN_121; // @[TLB.scala 252:34]
  wire  _GEN_122; // @[TLB.scala 252:34]
  wire  _GEN_123; // @[TLB.scala 249:72]
  wire  _GEN_124; // @[TLB.scala 249:72]
  wire  _GEN_125; // @[TLB.scala 249:72]
  wire  _GEN_126; // @[TLB.scala 249:72]
  wire  _T_1183; // @[TLB.scala 249:65]
  wire  _GEN_133; // @[TLB.scala 250:32]
  wire  _GEN_134; // @[TLB.scala 250:32]
  wire  _GEN_135; // @[TLB.scala 250:32]
  wire  _GEN_136; // @[TLB.scala 250:32]
  wire  _GEN_137; // @[TLB.scala 122:16]
  wire  _GEN_138; // @[TLB.scala 122:16]
  wire  _GEN_139; // @[TLB.scala 122:16]
  wire  _GEN_140; // @[TLB.scala 122:16]
  wire  _GEN_145; // @[TLB.scala 252:34]
  wire  _GEN_146; // @[TLB.scala 252:34]
  wire  _GEN_147; // @[TLB.scala 252:34]
  wire  _GEN_148; // @[TLB.scala 252:34]
  wire  _GEN_149; // @[TLB.scala 249:72]
  wire  _GEN_150; // @[TLB.scala 249:72]
  wire  _GEN_151; // @[TLB.scala 249:72]
  wire  _GEN_152; // @[TLB.scala 249:72]
  wire  _T_1201; // @[TLB.scala 249:65]
  wire  _GEN_159; // @[TLB.scala 250:32]
  wire  _GEN_160; // @[TLB.scala 250:32]
  wire  _GEN_161; // @[TLB.scala 250:32]
  wire  _GEN_162; // @[TLB.scala 250:32]
  wire  _GEN_163; // @[TLB.scala 122:16]
  wire  _GEN_164; // @[TLB.scala 122:16]
  wire  _GEN_165; // @[TLB.scala 122:16]
  wire  _GEN_166; // @[TLB.scala 122:16]
  wire  _GEN_171; // @[TLB.scala 252:34]
  wire  _GEN_172; // @[TLB.scala 252:34]
  wire  _GEN_173; // @[TLB.scala 252:34]
  wire  _GEN_174; // @[TLB.scala 252:34]
  wire  _GEN_175; // @[TLB.scala 249:72]
  wire  _GEN_176; // @[TLB.scala 249:72]
  wire  _GEN_177; // @[TLB.scala 249:72]
  wire  _GEN_178; // @[TLB.scala 249:72]
  wire  _T_1219; // @[TLB.scala 249:65]
  wire  _GEN_185; // @[TLB.scala 250:32]
  wire  _GEN_186; // @[TLB.scala 250:32]
  wire  _GEN_187; // @[TLB.scala 250:32]
  wire  _GEN_188; // @[TLB.scala 250:32]
  wire  _GEN_189; // @[TLB.scala 122:16]
  wire  _GEN_190; // @[TLB.scala 122:16]
  wire  _GEN_191; // @[TLB.scala 122:16]
  wire  _GEN_192; // @[TLB.scala 122:16]
  wire  _GEN_197; // @[TLB.scala 252:34]
  wire  _GEN_198; // @[TLB.scala 252:34]
  wire  _GEN_199; // @[TLB.scala 252:34]
  wire  _GEN_200; // @[TLB.scala 252:34]
  wire  _GEN_201; // @[TLB.scala 249:72]
  wire  _GEN_202; // @[TLB.scala 249:72]
  wire  _GEN_203; // @[TLB.scala 249:72]
  wire  _GEN_204; // @[TLB.scala 249:72]
  wire  _T_1237; // @[TLB.scala 249:65]
  wire  _GEN_211; // @[TLB.scala 250:32]
  wire  _GEN_212; // @[TLB.scala 250:32]
  wire  _GEN_213; // @[TLB.scala 250:32]
  wire  _GEN_214; // @[TLB.scala 250:32]
  wire  _GEN_215; // @[TLB.scala 122:16]
  wire  _GEN_216; // @[TLB.scala 122:16]
  wire  _GEN_217; // @[TLB.scala 122:16]
  wire  _GEN_218; // @[TLB.scala 122:16]
  wire  _GEN_223; // @[TLB.scala 252:34]
  wire  _GEN_224; // @[TLB.scala 252:34]
  wire  _GEN_225; // @[TLB.scala 252:34]
  wire  _GEN_226; // @[TLB.scala 252:34]
  wire  _GEN_227; // @[TLB.scala 249:72]
  wire  _GEN_228; // @[TLB.scala 249:72]
  wire  _GEN_229; // @[TLB.scala 249:72]
  wire  _GEN_230; // @[TLB.scala 249:72]
  wire  _T_1255; // @[TLB.scala 249:65]
  wire  _GEN_237; // @[TLB.scala 250:32]
  wire  _GEN_238; // @[TLB.scala 250:32]
  wire  _GEN_239; // @[TLB.scala 250:32]
  wire  _GEN_240; // @[TLB.scala 250:32]
  wire  _GEN_241; // @[TLB.scala 122:16]
  wire  _GEN_242; // @[TLB.scala 122:16]
  wire  _GEN_243; // @[TLB.scala 122:16]
  wire  _GEN_244; // @[TLB.scala 122:16]
  wire  _GEN_249; // @[TLB.scala 252:34]
  wire  _GEN_250; // @[TLB.scala 252:34]
  wire  _GEN_251; // @[TLB.scala 252:34]
  wire  _GEN_252; // @[TLB.scala 252:34]
  wire  _GEN_253; // @[TLB.scala 249:72]
  wire  _GEN_254; // @[TLB.scala 249:72]
  wire  _GEN_255; // @[TLB.scala 249:72]
  wire  _GEN_256; // @[TLB.scala 249:72]
  wire  _T_1273; // @[TLB.scala 249:65]
  wire  _GEN_263; // @[TLB.scala 250:32]
  wire  _GEN_264; // @[TLB.scala 250:32]
  wire  _GEN_265; // @[TLB.scala 250:32]
  wire  _GEN_266; // @[TLB.scala 250:32]
  wire  _GEN_267; // @[TLB.scala 122:16]
  wire  _GEN_268; // @[TLB.scala 122:16]
  wire  _GEN_269; // @[TLB.scala 122:16]
  wire  _GEN_270; // @[TLB.scala 122:16]
  wire  _GEN_275; // @[TLB.scala 252:34]
  wire  _GEN_276; // @[TLB.scala 252:34]
  wire  _GEN_277; // @[TLB.scala 252:34]
  wire  _GEN_278; // @[TLB.scala 252:34]
  wire  _GEN_279; // @[TLB.scala 249:72]
  wire  _GEN_280; // @[TLB.scala 249:72]
  wire  _GEN_281; // @[TLB.scala 249:72]
  wire  _GEN_282; // @[TLB.scala 249:72]
  wire  _GEN_291; // @[TLB.scala 242:54]
  wire  _GEN_295; // @[TLB.scala 242:54]
  wire  _GEN_299; // @[TLB.scala 242:54]
  wire  _GEN_303; // @[TLB.scala 242:54]
  wire  _GEN_305; // @[TLB.scala 242:54]
  wire  _GEN_306; // @[TLB.scala 242:54]
  wire  _GEN_307; // @[TLB.scala 242:54]
  wire  _GEN_308; // @[TLB.scala 242:54]
  wire  _GEN_315; // @[TLB.scala 242:54]
  wire  _GEN_316; // @[TLB.scala 242:54]
  wire  _GEN_317; // @[TLB.scala 242:54]
  wire  _GEN_318; // @[TLB.scala 242:54]
  wire  _GEN_325; // @[TLB.scala 242:54]
  wire  _GEN_326; // @[TLB.scala 242:54]
  wire  _GEN_327; // @[TLB.scala 242:54]
  wire  _GEN_328; // @[TLB.scala 242:54]
  wire  _GEN_335; // @[TLB.scala 242:54]
  wire  _GEN_336; // @[TLB.scala 242:54]
  wire  _GEN_337; // @[TLB.scala 242:54]
  wire  _GEN_338; // @[TLB.scala 242:54]
  wire  _GEN_345; // @[TLB.scala 242:54]
  wire  _GEN_346; // @[TLB.scala 242:54]
  wire  _GEN_347; // @[TLB.scala 242:54]
  wire  _GEN_348; // @[TLB.scala 242:54]
  wire  _GEN_355; // @[TLB.scala 242:54]
  wire  _GEN_356; // @[TLB.scala 242:54]
  wire  _GEN_357; // @[TLB.scala 242:54]
  wire  _GEN_358; // @[TLB.scala 242:54]
  wire  _GEN_365; // @[TLB.scala 242:54]
  wire  _GEN_366; // @[TLB.scala 242:54]
  wire  _GEN_367; // @[TLB.scala 242:54]
  wire  _GEN_368; // @[TLB.scala 242:54]
  wire  _GEN_375; // @[TLB.scala 242:54]
  wire  _GEN_376; // @[TLB.scala 242:54]
  wire  _GEN_377; // @[TLB.scala 242:54]
  wire  _GEN_378; // @[TLB.scala 242:54]
  wire  _GEN_387; // @[TLB.scala 237:68]
  wire  _GEN_391; // @[TLB.scala 237:68]
  wire  _GEN_395; // @[TLB.scala 237:68]
  wire  _GEN_399; // @[TLB.scala 237:68]
  wire  _GEN_403; // @[TLB.scala 237:68]
  wire  _GEN_405; // @[TLB.scala 237:68]
  wire  _GEN_406; // @[TLB.scala 237:68]
  wire  _GEN_407; // @[TLB.scala 237:68]
  wire  _GEN_408; // @[TLB.scala 237:68]
  wire  _GEN_415; // @[TLB.scala 237:68]
  wire  _GEN_416; // @[TLB.scala 237:68]
  wire  _GEN_417; // @[TLB.scala 237:68]
  wire  _GEN_418; // @[TLB.scala 237:68]
  wire  _GEN_425; // @[TLB.scala 237:68]
  wire  _GEN_426; // @[TLB.scala 237:68]
  wire  _GEN_427; // @[TLB.scala 237:68]
  wire  _GEN_428; // @[TLB.scala 237:68]
  wire  _GEN_435; // @[TLB.scala 237:68]
  wire  _GEN_436; // @[TLB.scala 237:68]
  wire  _GEN_437; // @[TLB.scala 237:68]
  wire  _GEN_438; // @[TLB.scala 237:68]
  wire  _GEN_445; // @[TLB.scala 237:68]
  wire  _GEN_446; // @[TLB.scala 237:68]
  wire  _GEN_447; // @[TLB.scala 237:68]
  wire  _GEN_448; // @[TLB.scala 237:68]
  wire  _GEN_455; // @[TLB.scala 237:68]
  wire  _GEN_456; // @[TLB.scala 237:68]
  wire  _GEN_457; // @[TLB.scala 237:68]
  wire  _GEN_458; // @[TLB.scala 237:68]
  wire  _GEN_465; // @[TLB.scala 237:68]
  wire  _GEN_466; // @[TLB.scala 237:68]
  wire  _GEN_467; // @[TLB.scala 237:68]
  wire  _GEN_468; // @[TLB.scala 237:68]
  wire  _GEN_475; // @[TLB.scala 237:68]
  wire  _GEN_476; // @[TLB.scala 237:68]
  wire  _GEN_477; // @[TLB.scala 237:68]
  wire  _GEN_478; // @[TLB.scala 237:68]
  wire  _GEN_487; // @[TLB.scala 217:20]
  wire  _GEN_491; // @[TLB.scala 217:20]
  wire  _GEN_495; // @[TLB.scala 217:20]
  wire  _GEN_499; // @[TLB.scala 217:20]
  wire  _GEN_503; // @[TLB.scala 217:20]
  wire  _GEN_505; // @[TLB.scala 217:20]
  wire  _GEN_506; // @[TLB.scala 217:20]
  wire  _GEN_507; // @[TLB.scala 217:20]
  wire  _GEN_508; // @[TLB.scala 217:20]
  wire  _GEN_515; // @[TLB.scala 217:20]
  wire  _GEN_516; // @[TLB.scala 217:20]
  wire  _GEN_517; // @[TLB.scala 217:20]
  wire  _GEN_518; // @[TLB.scala 217:20]
  wire  _GEN_525; // @[TLB.scala 217:20]
  wire  _GEN_526; // @[TLB.scala 217:20]
  wire  _GEN_527; // @[TLB.scala 217:20]
  wire  _GEN_528; // @[TLB.scala 217:20]
  wire  _GEN_535; // @[TLB.scala 217:20]
  wire  _GEN_536; // @[TLB.scala 217:20]
  wire  _GEN_537; // @[TLB.scala 217:20]
  wire  _GEN_538; // @[TLB.scala 217:20]
  wire  _GEN_545; // @[TLB.scala 217:20]
  wire  _GEN_546; // @[TLB.scala 217:20]
  wire  _GEN_547; // @[TLB.scala 217:20]
  wire  _GEN_548; // @[TLB.scala 217:20]
  wire  _GEN_555; // @[TLB.scala 217:20]
  wire  _GEN_556; // @[TLB.scala 217:20]
  wire  _GEN_557; // @[TLB.scala 217:20]
  wire  _GEN_558; // @[TLB.scala 217:20]
  wire  _GEN_565; // @[TLB.scala 217:20]
  wire  _GEN_566; // @[TLB.scala 217:20]
  wire  _GEN_567; // @[TLB.scala 217:20]
  wire  _GEN_568; // @[TLB.scala 217:20]
  wire  _GEN_575; // @[TLB.scala 217:20]
  wire  _GEN_576; // @[TLB.scala 217:20]
  wire  _GEN_577; // @[TLB.scala 217:20]
  wire  _GEN_578; // @[TLB.scala 217:20]
  wire [5:0] _T_1761; // @[Cat.scala 29:58]
  wire [13:0] ptw_ae_array; // @[Cat.scala 29:58]
  wire  _T_1770; // @[TLB.scala 261:32]
  wire [5:0] _T_1775; // @[Cat.scala 29:58]
  wire [12:0] _T_1782; // @[Cat.scala 29:58]
  wire [12:0] _T_1783; // @[TLB.scala 261:23]
  wire [12:0] _T_1797; // @[TLB.scala 261:89]
  wire [12:0] priv_rw_ok; // @[TLB.scala 261:84]
  wire [5:0] _T_1827; // @[Cat.scala 29:58]
  wire [12:0] _T_1834; // @[Cat.scala 29:58]
  wire [5:0] _T_1839; // @[Cat.scala 29:58]
  wire [12:0] _T_1846; // @[Cat.scala 29:58]
  wire [12:0] _T_1847; // @[TLB.scala 263:73]
  wire [12:0] _T_1848; // @[TLB.scala 263:68]
  wire [12:0] _T_1849; // @[TLB.scala 263:40]
  wire [13:0] r_array; // @[Cat.scala 29:58]
  wire [5:0] _T_1854; // @[Cat.scala 29:58]
  wire [12:0] _T_1861; // @[Cat.scala 29:58]
  wire [12:0] _T_1862; // @[TLB.scala 264:40]
  wire [13:0] w_array; // @[Cat.scala 29:58]
  wire [1:0] _T_1877; // @[Bitwise.scala 72:12]
  wire [5:0] _T_1882; // @[Cat.scala 29:58]
  wire [13:0] _T_1889; // @[Cat.scala 29:58]
  wire [13:0] pr_array; // @[TLB.scala 266:87]
  wire [1:0] _T_1892; // @[Bitwise.scala 72:12]
  wire [5:0] _T_1897; // @[Cat.scala 29:58]
  wire [13:0] _T_1904; // @[Cat.scala 29:58]
  wire [13:0] pw_array; // @[TLB.scala 267:87]
  wire [1:0] _T_1922; // @[Bitwise.scala 72:12]
  wire [5:0] _T_1927; // @[Cat.scala 29:58]
  wire [13:0] eff_array; // @[Cat.scala 29:58]
  wire [1:0] _T_1935; // @[Bitwise.scala 72:12]
  wire [5:0] _T_1940; // @[Cat.scala 29:58]
  wire [13:0] c_array; // @[Cat.scala 29:58]
  wire [1:0] _T_1948; // @[Bitwise.scala 72:12]
  wire [5:0] _T_1953; // @[Cat.scala 29:58]
  wire [13:0] ppp_array; // @[Cat.scala 29:58]
  wire [1:0] _T_1961; // @[Bitwise.scala 72:12]
  wire [5:0] _T_1966; // @[Cat.scala 29:58]
  wire [13:0] paa_array; // @[Cat.scala 29:58]
  wire [5:0] _T_1979; // @[Cat.scala 29:58]
  wire [13:0] pal_array; // @[Cat.scala 29:58]
  wire [13:0] ppp_array_if_cached; // @[TLB.scala 274:39]
  wire [13:0] paa_array_if_cached; // @[TLB.scala 275:39]
  wire [13:0] pal_array_if_cached; // @[TLB.scala 276:39]
  wire [3:0] _T_2001; // @[OneHot.scala 58:35]
  wire [3:0] _T_2003; // @[TLB.scala 279:69]
  wire [39:0] _GEN_1027; // @[TLB.scala 279:39]
  wire [39:0] _T_2004; // @[TLB.scala 279:39]
  wire  misaligned; // @[TLB.scala 279:75]
  wire [39:0] _T_2005; // @[TLB.scala 285:43]
  wire  _T_2007; // @[TLB.scala 286:61]
  wire  _T_2008; // @[TLB.scala 286:82]
  wire  _T_2009; // @[TLB.scala 286:67]
  wire  bad_va; // @[TLB.scala 280:117]
  wire  _T_2012; // @[package.scala 15:47]
  wire  _T_2013; // @[package.scala 15:47]
  wire  cmd_lrsc; // @[package.scala 64:59]
  wire  _T_2015; // @[package.scala 15:47]
  wire  _T_2016; // @[package.scala 15:47]
  wire  _T_2017; // @[package.scala 15:47]
  wire  _T_2018; // @[package.scala 15:47]
  wire  _T_2019; // @[package.scala 64:59]
  wire  _T_2020; // @[package.scala 64:59]
  wire  cmd_amo_logical; // @[package.scala 64:59]
  wire  _T_2022; // @[package.scala 15:47]
  wire  _T_2023; // @[package.scala 15:47]
  wire  _T_2024; // @[package.scala 15:47]
  wire  _T_2025; // @[package.scala 15:47]
  wire  _T_2026; // @[package.scala 15:47]
  wire  _T_2027; // @[package.scala 64:59]
  wire  _T_2028; // @[package.scala 64:59]
  wire  _T_2029; // @[package.scala 64:59]
  wire  cmd_amo_arithmetic; // @[package.scala 64:59]
  wire  cmd_put_partial; // @[TLB.scala 293:41]
  wire  _T_2031; // @[Consts.scala 82:31]
  wire  _T_2033; // @[Consts.scala 82:41]
  wire  _T_2035; // @[Consts.scala 82:58]
  wire  _T_2052; // @[Consts.scala 80:44]
  wire  cmd_read; // @[Consts.scala 82:75]
  wire  _T_2053; // @[Consts.scala 83:32]
  wire  _T_2055; // @[Consts.scala 83:42]
  wire  _T_2057; // @[Consts.scala 83:59]
  wire  cmd_write; // @[Consts.scala 83:76]
  wire  _T_2075; // @[package.scala 15:47]
  wire  _T_2076; // @[package.scala 15:47]
  wire  _T_2077; // @[package.scala 64:59]
  wire  cmd_write_perms; // @[TLB.scala 296:35]
  wire [13:0] _T_2078; // @[TLB.scala 301:8]
  wire [13:0] _T_2080; // @[TLB.scala 302:8]
  wire [13:0] ae_array; // @[TLB.scala 301:37]
  wire [13:0] _T_2082; // @[TLB.scala 303:44]
  wire [13:0] ae_ld_array; // @[TLB.scala 303:24]
  wire [13:0] _T_2084; // @[TLB.scala 305:35]
  wire [13:0] _T_2085; // @[TLB.scala 305:8]
  wire [13:0] _T_2087; // @[TLB.scala 306:8]
  wire [13:0] _T_2088; // @[TLB.scala 305:53]
  wire [13:0] _T_2090; // @[TLB.scala 307:8]
  wire [13:0] _T_2091; // @[TLB.scala 306:53]
  wire [13:0] _T_2093; // @[TLB.scala 308:8]
  wire [13:0] ae_st_array; // @[TLB.scala 307:53]
  wire  _T_2104; // @[TLB.scala 314:36]
  wire [13:0] ma_ld_array; // @[TLB.scala 314:24]
  wire  _T_2106; // @[TLB.scala 315:36]
  wire [13:0] ma_st_array; // @[TLB.scala 315:24]
  wire [13:0] _T_2108; // @[TLB.scala 316:45]
  wire [13:0] pf_ld_array; // @[TLB.scala 316:24]
  wire [13:0] _T_2110; // @[TLB.scala 317:52]
  wire [13:0] pf_st_array; // @[TLB.scala 317:24]
  wire  tlb_hit; // @[TLB.scala 320:27]
  wire  _T_2114; // @[TLB.scala 321:29]
  wire  tlb_miss; // @[TLB.scala 321:40]
  reg [6:0] _T_2116; // @[Replacement.scala 158:30]
  reg [31:0] _RAND_98;
  reg [2:0] _T_2117; // @[Replacement.scala 158:30]
  reg [31:0] _RAND_99;
  wire  _T_2118; // @[TLB.scala 325:22]
  wire  _T_2119; // @[package.scala 64:59]
  wire  _T_2120; // @[package.scala 64:59]
  wire  _T_2121; // @[package.scala 64:59]
  wire  _T_2122; // @[package.scala 64:59]
  wire  _T_2123; // @[package.scala 64:59]
  wire  _T_2124; // @[package.scala 64:59]
  wire  _T_2125; // @[package.scala 64:59]
  wire [7:0] _T_2132; // @[Cat.scala 29:58]
  wire  _T_2135; // @[OneHot.scala 32:14]
  wire [3:0] _T_2136; // @[OneHot.scala 32:28]
  wire  _T_2139; // @[OneHot.scala 32:14]
  wire [1:0] _T_2140; // @[OneHot.scala 32:28]
  wire [2:0] _T_2143; // @[Cat.scala 29:58]
  wire  _T_2157; // @[Replacement.scala 193:16]
  wire  _T_2161; // @[Replacement.scala 196:16]
  wire [2:0] _T_2163; // @[Cat.scala 29:58]
  wire [2:0] _T_2164; // @[Replacement.scala 193:16]
  wire  _T_2173; // @[Replacement.scala 193:16]
  wire  _T_2177; // @[Replacement.scala 196:16]
  wire [2:0] _T_2179; // @[Cat.scala 29:58]
  wire [2:0] _T_2180; // @[Replacement.scala 196:16]
  wire [6:0] _T_2182; // @[Cat.scala 29:58]
  wire  _T_2183; // @[package.scala 64:59]
  wire  _T_2184; // @[package.scala 64:59]
  wire  _T_2185; // @[package.scala 64:59]
  wire [3:0] _T_2188; // @[Cat.scala 29:58]
  wire  _T_2191; // @[OneHot.scala 32:14]
  wire [1:0] _T_2192; // @[OneHot.scala 32:28]
  wire [1:0] _T_2194; // @[Cat.scala 29:58]
  wire  _T_2203; // @[Replacement.scala 193:16]
  wire  _T_2207; // @[Replacement.scala 196:16]
  wire [2:0] _T_2209; // @[Cat.scala 29:58]
  wire  _T_2219; // @[Misc.scala 182:16]
  wire  _T_2221; // @[Misc.scala 182:61]
  wire  _T_2223; // @[Misc.scala 182:16]
  wire  _T_2225; // @[Misc.scala 182:61]
  wire  _T_2226; // @[Misc.scala 182:49]
  wire  _T_2235; // @[Misc.scala 182:16]
  wire  _T_2237; // @[Misc.scala 182:61]
  wire  _T_2239; // @[Misc.scala 182:16]
  wire  _T_2241; // @[Misc.scala 182:61]
  wire  _T_2242; // @[Misc.scala 182:49]
  wire  _T_2243; // @[Misc.scala 182:16]
  wire  _T_2244; // @[Misc.scala 182:37]
  wire  _T_2245; // @[Misc.scala 182:61]
  wire  _T_2246; // @[Misc.scala 182:49]
  wire  _T_2256; // @[Misc.scala 182:16]
  wire  _T_2258; // @[Misc.scala 182:61]
  wire  _T_2260; // @[Misc.scala 182:16]
  wire  _T_2262; // @[Misc.scala 182:61]
  wire  _T_2263; // @[Misc.scala 182:49]
  wire  _T_2270; // @[Misc.scala 182:16]
  wire  _T_2272; // @[Misc.scala 182:61]
  wire  _T_2279; // @[Misc.scala 182:16]
  wire  _T_2281; // @[Misc.scala 182:61]
  wire  _T_2283; // @[Misc.scala 182:16]
  wire  _T_2284; // @[Misc.scala 182:37]
  wire  _T_2285; // @[Misc.scala 182:61]
  wire  _T_2286; // @[Misc.scala 182:49]
  wire  _T_2287; // @[Misc.scala 182:16]
  wire  _T_2288; // @[Misc.scala 182:37]
  wire  _T_2289; // @[Misc.scala 182:61]
  wire  _T_2290; // @[Misc.scala 182:49]
  wire  _T_2292; // @[Misc.scala 182:37]
  wire  _T_2293; // @[Misc.scala 182:61]
  wire  multipleHits; // @[Misc.scala 182:49]
  wire  _T_2295; // @[TLB.scala 338:28]
  wire [13:0] _T_2296; // @[TLB.scala 338:57]
  wire  _T_2297; // @[TLB.scala 338:65]
  wire  _T_2299; // @[TLB.scala 339:28]
  wire [13:0] _T_2300; // @[TLB.scala 339:64]
  wire  _T_2301; // @[TLB.scala 339:72]
  wire [13:0] _T_2306; // @[TLB.scala 341:33]
  wire [13:0] _T_2308; // @[TLB.scala 342:33]
  wire [13:0] _T_2313; // @[TLB.scala 344:33]
  wire [13:0] _T_2315; // @[TLB.scala 345:33]
  wire [13:0] _T_2317; // @[TLB.scala 347:33]
  wire  _T_2324; // @[TLB.scala 350:29]
  wire  _T_2330; // @[Decoupled.scala 40:37]
  wire  _T_2331; // @[TLB.scala 359:25]
  wire  _T_2337; // @[Replacement.scala 240:16]
  wire [1:0] _T_2338; // @[Cat.scala 29:58]
  wire [3:0] _T_2341; // @[Cat.scala 29:58]
  wire  _T_2342; // @[TLB.scala 407:16]
  wire  _T_2344; // @[OneHot.scala 47:40]
  wire  _T_2345; // @[OneHot.scala 47:40]
  wire  _T_2346; // @[OneHot.scala 47:40]
  wire  _T_2360; // @[Replacement.scala 240:16]
  wire [1:0] _T_2361; // @[Cat.scala 29:58]
  wire  _T_2367; // @[Replacement.scala 240:16]
  wire [1:0] _T_2368; // @[Cat.scala 29:58]
  wire [1:0] _T_2369; // @[Replacement.scala 240:16]
  wire [2:0] _T_2370; // @[Cat.scala 29:58]
  wire [7:0] _T_2401; // @[Cat.scala 29:58]
  wire  _T_2402; // @[TLB.scala 407:16]
  wire  _T_2404; // @[OneHot.scala 47:40]
  wire  _T_2405; // @[OneHot.scala 47:40]
  wire  _T_2406; // @[OneHot.scala 47:40]
  wire  _T_2407; // @[OneHot.scala 47:40]
  wire  _T_2408; // @[OneHot.scala 47:40]
  wire  _T_2409; // @[OneHot.scala 47:40]
  wire  _T_2410; // @[OneHot.scala 47:40]
  wire  _T_2447; // @[TLB.scala 373:17]
  wire  _T_2448; // @[TLB.scala 373:28]
  wire  _T_2451; // @[TLB.scala 381:72]
  wire  _T_2452; // @[TLB.scala 381:34]
  wire  _T_2454; // @[TLB.scala 381:13]
  wire  _T_2462; // @[TLB.scala 135:61]
  wire  _GEN_681; // @[TLB.scala 143:19]
  wire  _GEN_682; // @[TLB.scala 143:19]
  wire  _GEN_683; // @[TLB.scala 143:19]
  wire  _GEN_684; // @[TLB.scala 143:19]
  wire  _GEN_685; // @[TLB.scala 384:40]
  wire  _GEN_686; // @[TLB.scala 384:40]
  wire  _GEN_687; // @[TLB.scala 384:40]
  wire  _GEN_688; // @[TLB.scala 384:40]
  wire  _T_2617; // @[TLB.scala 135:61]
  wire  _GEN_709; // @[TLB.scala 143:19]
  wire  _GEN_710; // @[TLB.scala 143:19]
  wire  _GEN_711; // @[TLB.scala 143:19]
  wire  _GEN_712; // @[TLB.scala 143:19]
  wire  _GEN_713; // @[TLB.scala 384:40]
  wire  _GEN_714; // @[TLB.scala 384:40]
  wire  _GEN_715; // @[TLB.scala 384:40]
  wire  _GEN_716; // @[TLB.scala 384:40]
  wire  _T_2772; // @[TLB.scala 135:61]
  wire  _GEN_737; // @[TLB.scala 143:19]
  wire  _GEN_738; // @[TLB.scala 143:19]
  wire  _GEN_739; // @[TLB.scala 143:19]
  wire  _GEN_740; // @[TLB.scala 143:19]
  wire  _GEN_741; // @[TLB.scala 384:40]
  wire  _GEN_742; // @[TLB.scala 384:40]
  wire  _GEN_743; // @[TLB.scala 384:40]
  wire  _GEN_744; // @[TLB.scala 384:40]
  wire  _T_2927; // @[TLB.scala 135:61]
  wire  _GEN_765; // @[TLB.scala 143:19]
  wire  _GEN_766; // @[TLB.scala 143:19]
  wire  _GEN_767; // @[TLB.scala 143:19]
  wire  _GEN_768; // @[TLB.scala 143:19]
  wire  _GEN_769; // @[TLB.scala 384:40]
  wire  _GEN_770; // @[TLB.scala 384:40]
  wire  _GEN_771; // @[TLB.scala 384:40]
  wire  _GEN_772; // @[TLB.scala 384:40]
  wire  _T_3082; // @[TLB.scala 135:61]
  wire  _GEN_793; // @[TLB.scala 143:19]
  wire  _GEN_794; // @[TLB.scala 143:19]
  wire  _GEN_795; // @[TLB.scala 143:19]
  wire  _GEN_796; // @[TLB.scala 143:19]
  wire  _GEN_797; // @[TLB.scala 384:40]
  wire  _GEN_798; // @[TLB.scala 384:40]
  wire  _GEN_799; // @[TLB.scala 384:40]
  wire  _GEN_800; // @[TLB.scala 384:40]
  wire  _T_3237; // @[TLB.scala 135:61]
  wire  _GEN_821; // @[TLB.scala 143:19]
  wire  _GEN_822; // @[TLB.scala 143:19]
  wire  _GEN_823; // @[TLB.scala 143:19]
  wire  _GEN_824; // @[TLB.scala 143:19]
  wire  _GEN_825; // @[TLB.scala 384:40]
  wire  _GEN_826; // @[TLB.scala 384:40]
  wire  _GEN_827; // @[TLB.scala 384:40]
  wire  _GEN_828; // @[TLB.scala 384:40]
  wire  _T_3392; // @[TLB.scala 135:61]
  wire  _GEN_849; // @[TLB.scala 143:19]
  wire  _GEN_850; // @[TLB.scala 143:19]
  wire  _GEN_851; // @[TLB.scala 143:19]
  wire  _GEN_852; // @[TLB.scala 143:19]
  wire  _GEN_853; // @[TLB.scala 384:40]
  wire  _GEN_854; // @[TLB.scala 384:40]
  wire  _GEN_855; // @[TLB.scala 384:40]
  wire  _GEN_856; // @[TLB.scala 384:40]
  wire  _T_3547; // @[TLB.scala 135:61]
  wire  _GEN_877; // @[TLB.scala 143:19]
  wire  _GEN_878; // @[TLB.scala 143:19]
  wire  _GEN_879; // @[TLB.scala 143:19]
  wire  _GEN_880; // @[TLB.scala 143:19]
  wire  _GEN_881; // @[TLB.scala 384:40]
  wire  _GEN_882; // @[TLB.scala 384:40]
  wire  _GEN_883; // @[TLB.scala 384:40]
  wire  _GEN_884; // @[TLB.scala 384:40]
  wire  _GEN_890; // @[TLB.scala 143:19]
  wire  _GEN_891; // @[TLB.scala 384:40]
  wire  _GEN_894; // @[TLB.scala 143:19]
  wire  _GEN_895; // @[TLB.scala 384:40]
  wire  _GEN_898; // @[TLB.scala 143:19]
  wire  _GEN_899; // @[TLB.scala 384:40]
  wire  _GEN_902; // @[TLB.scala 143:19]
  wire  _GEN_903; // @[TLB.scala 384:40]
  wire  _GEN_906; // @[TLB.scala 143:19]
  wire  _GEN_907; // @[TLB.scala 384:40]
  wire  _T_3897; // @[TLB.scala 388:24]
  reg [19:0] TLB_state; // @[Register tracking TLB state]
  reg [31:0] _RAND_100;
  reg  TLB_cov [0:1048575]; // @[Coverage map for TLB]
  reg [31:0] _RAND_101;
  wire  TLB_cov_read_data; // @[Coverage map for TLB]
  wire [19:0] TLB_cov_read_addr; // @[Coverage map for TLB]
  wire  TLB_cov_write_data; // @[Coverage map for TLB]
  wire [19:0] TLB_cov_write_addr; // @[Coverage map for TLB]
  wire  TLB_cov_write_mask; // @[Coverage map for TLB]
  wire  TLB_cov_write_en; // @[Coverage map for TLB]
  reg [29:0] TLB_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_102;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire  mux_cond_6;
  wire  mux_cond_7;
  wire  mux_cond_8;
  wire  mux_cond_9;
  wire  mux_cond_10;
  wire  mux_cond_11;
  wire  mux_cond_12;
  wire  mux_cond_13;
  wire  mux_cond_14;
  wire  mux_cond_15;
  wire  mux_cond_16;
  wire  mux_cond_17;
  wire  mux_cond_18;
  wire  mux_cond_19;
  wire  mux_cond_20;
  wire  mux_cond_21;
  wire  mux_cond_22;
  wire  mux_cond_23;
  wire  mux_cond_24;
  wire  mux_cond_25;
  wire  mux_cond_26;
  wire  mux_cond_27;
  wire  mux_cond_28;
  wire  mux_cond_29;
  wire  mux_cond_30;
  wire  mux_cond_31;
  wire  mux_cond_32;
  wire  mux_cond_33;
  wire  mux_cond_34;
  wire  mux_cond_35;
  wire  mux_cond_36;
  wire  mux_cond_37;
  wire  mux_cond_38;
  wire  mux_cond_39;
  wire  mux_cond_40;
  wire  mux_cond_41;
  wire  mux_cond_42;
  wire  mux_cond_43;
  wire  mux_cond_44;
  wire  mux_cond_45;
  wire  mux_cond_46;
  wire  mux_cond_47;
  wire  mux_cond_48;
  wire  mux_cond_49;
  wire  mux_cond_50;
  wire  mux_cond_51;
  wire  mux_cond_52;
  wire  mux_cond_53;
  wire  mux_cond_54;
  wire  mux_cond_55;
  wire  mux_cond_56;
  wire  mux_cond_57;
  wire  mux_cond_58;
  wire  mux_cond_59;
  wire  mux_cond_60;
  wire  mux_cond_61;
  wire  mux_cond_62;
  wire  mux_cond_63;
  wire  mux_cond_64;
  wire  mux_cond_65;
  wire  mux_cond_66;
  wire  mux_cond_67;
  wire  mux_cond_68;
  wire [6:0] state_shl;
  wire [19:0] state_pad;
  wire [14:0] r_sectored_repl_addr_shl;
  wire [19:0] r_sectored_repl_addr_pad;
  wire [3:0] r_superpage_repl_addr_shl;
  wire [19:0] r_superpage_repl_addr_pad;
  wire [10:0] r_sectored_hit_addr_shl;
  wire [19:0] r_sectored_hit_addr_pad;
  wire [15:0] special_entry_valid_0_shl;
  wire [19:0] special_entry_valid_0_pad;
  wire [12:0] r_sectored_hit_shl;
  wire [19:0] r_sectored_hit_pad;
  wire [4:0] special_entry_level_shl;
  wire [19:0] special_entry_level_pad;
  wire [8:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [12:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [5:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [7:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [7:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [5:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [4:0] mux_cond_6_shl;
  wire [19:0] mux_cond_6_pad;
  wire [18:0] mux_cond_7_shl;
  wire [19:0] mux_cond_7_pad;
  wire [2:0] mux_cond_8_shl;
  wire [19:0] mux_cond_8_pad;
  wire [6:0] mux_cond_9_shl;
  wire [19:0] mux_cond_9_pad;
  wire  mux_cond_10_shl;
  wire [19:0] mux_cond_10_pad;
  wire [14:0] mux_cond_11_shl;
  wire [19:0] mux_cond_11_pad;
  wire [15:0] mux_cond_12_shl;
  wire [19:0] mux_cond_12_pad;
  wire  mux_cond_13_shl;
  wire [19:0] mux_cond_13_pad;
  wire [17:0] mux_cond_14_shl;
  wire [19:0] mux_cond_14_pad;
  wire [9:0] mux_cond_15_shl;
  wire [19:0] mux_cond_15_pad;
  wire [4:0] mux_cond_16_shl;
  wire [19:0] mux_cond_16_pad;
  wire [7:0] mux_cond_17_shl;
  wire [19:0] mux_cond_17_pad;
  wire [15:0] mux_cond_18_shl;
  wire [19:0] mux_cond_18_pad;
  wire [10:0] mux_cond_19_shl;
  wire [19:0] mux_cond_19_pad;
  wire [4:0] mux_cond_20_shl;
  wire [19:0] mux_cond_20_pad;
  wire [5:0] mux_cond_21_shl;
  wire [19:0] mux_cond_21_pad;
  wire [7:0] mux_cond_22_shl;
  wire [19:0] mux_cond_22_pad;
  wire [17:0] mux_cond_23_shl;
  wire [19:0] mux_cond_23_pad;
  wire [8:0] mux_cond_24_shl;
  wire [19:0] mux_cond_24_pad;
  wire [7:0] mux_cond_25_shl;
  wire [19:0] mux_cond_25_pad;
  wire [18:0] mux_cond_26_shl;
  wire [19:0] mux_cond_26_pad;
  wire [9:0] mux_cond_27_shl;
  wire [19:0] mux_cond_27_pad;
  wire [10:0] mux_cond_28_shl;
  wire [19:0] mux_cond_28_pad;
  wire [9:0] mux_cond_29_shl;
  wire [19:0] mux_cond_29_pad;
  wire [16:0] mux_cond_30_shl;
  wire [19:0] mux_cond_30_pad;
  wire [3:0] mux_cond_31_shl;
  wire [19:0] mux_cond_31_pad;
  wire [1:0] mux_cond_32_shl;
  wire [19:0] mux_cond_32_pad;
  wire [5:0] mux_cond_33_shl;
  wire [19:0] mux_cond_33_pad;
  wire [4:0] mux_cond_34_shl;
  wire [19:0] mux_cond_34_pad;
  wire [12:0] mux_cond_35_shl;
  wire [19:0] mux_cond_35_pad;
  wire [9:0] mux_cond_36_shl;
  wire [19:0] mux_cond_36_pad;
  wire [4:0] mux_cond_37_shl;
  wire [19:0] mux_cond_37_pad;
  wire [10:0] mux_cond_38_shl;
  wire [19:0] mux_cond_38_pad;
  wire [8:0] mux_cond_39_shl;
  wire [19:0] mux_cond_39_pad;
  wire [18:0] mux_cond_40_shl;
  wire [19:0] mux_cond_40_pad;
  wire [17:0] mux_cond_41_shl;
  wire [19:0] mux_cond_41_pad;
  wire [18:0] mux_cond_42_shl;
  wire [19:0] mux_cond_42_pad;
  wire [18:0] mux_cond_43_shl;
  wire [19:0] mux_cond_43_pad;
  wire  mux_cond_44_shl;
  wire [19:0] mux_cond_44_pad;
  wire [11:0] mux_cond_45_shl;
  wire [19:0] mux_cond_45_pad;
  wire [15:0] mux_cond_46_shl;
  wire [19:0] mux_cond_46_pad;
  wire [6:0] mux_cond_47_shl;
  wire [19:0] mux_cond_47_pad;
  wire  mux_cond_48_shl;
  wire [19:0] mux_cond_48_pad;
  wire [18:0] mux_cond_49_shl;
  wire [19:0] mux_cond_49_pad;
  wire [19:0] mux_cond_50_shl;
  wire [19:0] mux_cond_50_pad;
  wire [7:0] mux_cond_51_shl;
  wire [19:0] mux_cond_51_pad;
  wire [18:0] mux_cond_52_shl;
  wire [19:0] mux_cond_52_pad;
  wire [17:0] mux_cond_53_shl;
  wire [19:0] mux_cond_53_pad;
  wire [17:0] mux_cond_54_shl;
  wire [19:0] mux_cond_54_pad;
  wire [15:0] mux_cond_55_shl;
  wire [19:0] mux_cond_55_pad;
  wire [4:0] mux_cond_56_shl;
  wire [19:0] mux_cond_56_pad;
  wire [3:0] mux_cond_57_shl;
  wire [19:0] mux_cond_57_pad;
  wire [6:0] mux_cond_58_shl;
  wire [19:0] mux_cond_58_pad;
  wire [10:0] mux_cond_59_shl;
  wire [19:0] mux_cond_59_pad;
  wire [15:0] mux_cond_60_shl;
  wire [19:0] mux_cond_60_pad;
  wire [19:0] mux_cond_61_shl;
  wire [19:0] mux_cond_61_pad;
  wire [14:0] mux_cond_62_shl;
  wire [19:0] mux_cond_62_pad;
  wire [11:0] mux_cond_63_shl;
  wire [19:0] mux_cond_63_pad;
  wire [2:0] mux_cond_64_shl;
  wire [19:0] mux_cond_64_pad;
  wire [7:0] mux_cond_65_shl;
  wire [19:0] mux_cond_65_pad;
  wire [3:0] mux_cond_66_shl;
  wire [19:0] mux_cond_66_pad;
  wire [1:0] mux_cond_67_shl;
  wire [19:0] mux_cond_67_pad;
  wire [7:0] mux_cond_68_shl;
  wire [19:0] mux_cond_68_pad;
  wire [19:0] superpage_entries_2_level_shl;
  wire [19:0] superpage_entries_2_level_pad;
  wire [2:0] sectored_entries_7_valid_3_shl;
  wire [19:0] sectored_entries_7_valid_3_pad;
  wire [19:0] superpage_entries_1_level_shl;
  wire [19:0] superpage_entries_1_level_pad;
  wire [18:0] superpage_entries_1_valid_0_shl;
  wire [19:0] superpage_entries_1_valid_0_pad;
  wire [10:0] sectored_entries_3_valid_0_shl;
  wire [19:0] sectored_entries_3_valid_0_pad;
  wire [2:0] sectored_entries_1_valid_3_shl;
  wire [19:0] sectored_entries_1_valid_3_pad;
  wire [2:0] sectored_entries_6_valid_3_shl;
  wire [19:0] sectored_entries_6_valid_3_pad;
  wire [10:0] sectored_entries_1_valid_0_shl;
  wire [19:0] sectored_entries_1_valid_0_pad;
  wire [10:0] sectored_entries_2_valid_0_shl;
  wire [19:0] sectored_entries_2_valid_0_pad;
  wire [5:0] sectored_entries_3_valid_1_shl;
  wire [19:0] sectored_entries_3_valid_1_pad;
  wire [2:0] sectored_entries_5_valid_3_shl;
  wire [19:0] sectored_entries_5_valid_3_pad;
  wire [18:0] superpage_entries_3_valid_0_shl;
  wire [19:0] superpage_entries_3_valid_0_pad;
  wire [5:0] sectored_entries_5_valid_1_shl;
  wire [19:0] sectored_entries_5_valid_1_pad;
  wire [2:0] sectored_entries_0_valid_3_shl;
  wire [19:0] sectored_entries_0_valid_3_pad;
  wire [10:0] sectored_entries_6_valid_0_shl;
  wire [19:0] sectored_entries_6_valid_0_pad;
  wire [10:0] sectored_entries_0_valid_0_shl;
  wire [19:0] sectored_entries_0_valid_0_pad;
  wire [5:0] sectored_entries_4_valid_2_shl;
  wire [19:0] sectored_entries_4_valid_2_pad;
  wire [18:0] superpage_entries_2_valid_0_shl;
  wire [19:0] superpage_entries_2_valid_0_pad;
  wire [5:0] sectored_entries_2_valid_1_shl;
  wire [19:0] sectored_entries_2_valid_1_pad;
  wire [19:0] superpage_entries_0_level_shl;
  wire [19:0] superpage_entries_0_level_pad;
  wire [5:0] sectored_entries_1_valid_1_shl;
  wire [19:0] sectored_entries_1_valid_1_pad;
  wire [2:0] sectored_entries_4_valid_3_shl;
  wire [19:0] sectored_entries_4_valid_3_pad;
  wire [5:0] sectored_entries_0_valid_1_shl;
  wire [19:0] sectored_entries_0_valid_1_pad;
  wire [10:0] sectored_entries_4_valid_0_shl;
  wire [19:0] sectored_entries_4_valid_0_pad;
  wire [5:0] sectored_entries_0_valid_2_shl;
  wire [19:0] sectored_entries_0_valid_2_pad;
  wire [5:0] sectored_entries_1_valid_2_shl;
  wire [19:0] sectored_entries_1_valid_2_pad;
  wire [5:0] sectored_entries_2_valid_2_shl;
  wire [19:0] sectored_entries_2_valid_2_pad;
  wire [10:0] sectored_entries_7_valid_0_shl;
  wire [19:0] sectored_entries_7_valid_0_pad;
  wire [5:0] sectored_entries_5_valid_2_shl;
  wire [19:0] sectored_entries_5_valid_2_pad;
  wire [5:0] sectored_entries_7_valid_2_shl;
  wire [19:0] sectored_entries_7_valid_2_pad;
  wire [5:0] sectored_entries_4_valid_1_shl;
  wire [19:0] sectored_entries_4_valid_1_pad;
  wire [10:0] sectored_entries_5_valid_0_shl;
  wire [19:0] sectored_entries_5_valid_0_pad;
  wire [5:0] sectored_entries_7_valid_1_shl;
  wire [19:0] sectored_entries_7_valid_1_pad;
  wire [19:0] superpage_entries_3_level_shl;
  wire [19:0] superpage_entries_3_level_pad;
  wire [2:0] sectored_entries_3_valid_3_shl;
  wire [19:0] sectored_entries_3_valid_3_pad;
  wire [2:0] sectored_entries_2_valid_3_shl;
  wire [19:0] sectored_entries_2_valid_3_pad;
  wire [18:0] superpage_entries_0_valid_0_shl;
  wire [19:0] superpage_entries_0_valid_0_pad;
  wire [5:0] sectored_entries_6_valid_1_shl;
  wire [19:0] sectored_entries_6_valid_1_pad;
  wire [5:0] sectored_entries_3_valid_2_shl;
  wire [19:0] sectored_entries_3_valid_2_pad;
  wire [5:0] sectored_entries_6_valid_2_shl;
  wire [19:0] sectored_entries_6_valid_2_pad;
  wire [19:0] TLB_xor64;
  wire [19:0] TLB_xor31;
  wire [19:0] TLB_xor65;
  wire [19:0] TLB_xor66;
  wire [19:0] TLB_xor32;
  wire [19:0] TLB_xor15;
  wire [19:0] TLB_xor68;
  wire [19:0] TLB_xor33;
  wire [19:0] TLB_xor69;
  wire [19:0] TLB_xor70;
  wire [19:0] TLB_xor34;
  wire [19:0] TLB_xor16;
  wire [19:0] TLB_xor7;
  wire [19:0] TLB_xor72;
  wire [19:0] TLB_xor35;
  wire [19:0] TLB_xor73;
  wire [19:0] TLB_xor74;
  wire [19:0] TLB_xor36;
  wire [19:0] TLB_xor17;
  wire [19:0] TLB_xor75;
  wire [19:0] TLB_xor76;
  wire [19:0] TLB_xor37;
  wire [19:0] TLB_xor77;
  wire [19:0] TLB_xor78;
  wire [19:0] TLB_xor38;
  wire [19:0] TLB_xor18;
  wire [19:0] TLB_xor8;
  wire [19:0] TLB_xor3;
  wire [19:0] TLB_xor80;
  wire [19:0] TLB_xor39;
  wire [19:0] TLB_xor81;
  wire [19:0] TLB_xor82;
  wire [19:0] TLB_xor40;
  wire [19:0] TLB_xor19;
  wire [19:0] TLB_xor84;
  wire [19:0] TLB_xor41;
  wire [19:0] TLB_xor85;
  wire [19:0] TLB_xor86;
  wire [19:0] TLB_xor42;
  wire [19:0] TLB_xor20;
  wire [19:0] TLB_xor9;
  wire [19:0] TLB_xor88;
  wire [19:0] TLB_xor43;
  wire [19:0] TLB_xor89;
  wire [19:0] TLB_xor90;
  wire [19:0] TLB_xor44;
  wire [19:0] TLB_xor21;
  wire [19:0] TLB_xor91;
  wire [19:0] TLB_xor92;
  wire [19:0] TLB_xor45;
  wire [19:0] TLB_xor93;
  wire [19:0] TLB_xor94;
  wire [19:0] TLB_xor46;
  wire [19:0] TLB_xor22;
  wire [19:0] TLB_xor10;
  wire [19:0] TLB_xor4;
  wire [19:0] TLB_xor1;
  wire [19:0] TLB_xor96;
  wire [19:0] TLB_xor47;
  wire [19:0] TLB_xor97;
  wire [19:0] TLB_xor98;
  wire [19:0] TLB_xor48;
  wire [19:0] TLB_xor23;
  wire [19:0] TLB_xor100;
  wire [19:0] TLB_xor49;
  wire [19:0] TLB_xor101;
  wire [19:0] TLB_xor102;
  wire [19:0] TLB_xor50;
  wire [19:0] TLB_xor24;
  wire [19:0] TLB_xor11;
  wire [19:0] TLB_xor104;
  wire [19:0] TLB_xor51;
  wire [19:0] TLB_xor105;
  wire [19:0] TLB_xor106;
  wire [19:0] TLB_xor52;
  wire [19:0] TLB_xor25;
  wire [19:0] TLB_xor107;
  wire [19:0] TLB_xor108;
  wire [19:0] TLB_xor53;
  wire [19:0] TLB_xor109;
  wire [19:0] TLB_xor110;
  wire [19:0] TLB_xor54;
  wire [19:0] TLB_xor26;
  wire [19:0] TLB_xor12;
  wire [19:0] TLB_xor5;
  wire [19:0] TLB_xor112;
  wire [19:0] TLB_xor55;
  wire [19:0] TLB_xor113;
  wire [19:0] TLB_xor114;
  wire [19:0] TLB_xor56;
  wire [19:0] TLB_xor27;
  wire [19:0] TLB_xor116;
  wire [19:0] TLB_xor57;
  wire [19:0] TLB_xor117;
  wire [19:0] TLB_xor118;
  wire [19:0] TLB_xor58;
  wire [19:0] TLB_xor28;
  wire [19:0] TLB_xor13;
  wire [19:0] TLB_xor120;
  wire [19:0] TLB_xor59;
  wire [19:0] TLB_xor121;
  wire [19:0] TLB_xor122;
  wire [19:0] TLB_xor60;
  wire [19:0] TLB_xor29;
  wire [19:0] TLB_xor123;
  wire [19:0] TLB_xor124;
  wire [19:0] TLB_xor61;
  wire [19:0] TLB_xor125;
  wire [19:0] TLB_xor126;
  wire [19:0] TLB_xor62;
  wire [19:0] TLB_xor30;
  wire [19:0] TLB_xor14;
  wire [19:0] TLB_xor6;
  wire [19:0] TLB_xor2;
  wire [19:0] TLB_xor0;
  wire [29:0] OptimizationBarrier_20_sum;
  wire [29:0] OptimizationBarrier_21_sum;
  wire [29:0] OptimizationBarrier_35_sum;
  wire [29:0] OptimizationBarrier_6_sum;
  wire [29:0] OptimizationBarrier_16_sum;
  wire [29:0] OptimizationBarrier_12_sum;
  wire [29:0] OptimizationBarrier_9_sum;
  wire [29:0] OptimizationBarrier_8_sum;
  wire [29:0] OptimizationBarrier_2_sum;
  wire [29:0] OptimizationBarrier_25_sum;
  wire [29:0] pmp_sum;
  wire [29:0] OptimizationBarrier_23_sum;
  wire [29:0] OptimizationBarrier_27_sum;
  wire [29:0] OptimizationBarrier_30_sum;
  wire [29:0] OptimizationBarrier_1_sum;
  wire [29:0] OptimizationBarrier_18_sum;
  wire [29:0] OptimizationBarrier_31_sum;
  wire [29:0] OptimizationBarrier_19_sum;
  wire [29:0] OptimizationBarrier_37_sum;
  wire [29:0] OptimizationBarrier_28_sum;
  wire [29:0] OptimizationBarrier_33_sum;
  wire [29:0] OptimizationBarrier_4_sum;
  wire [29:0] OptimizationBarrier_38_sum;
  wire [29:0] OptimizationBarrier_sum;
  wire [29:0] OptimizationBarrier_34_sum;
  wire [29:0] OptimizationBarrier_24_sum;
  wire [29:0] OptimizationBarrier_22_sum;
  wire [29:0] OptimizationBarrier_10_sum;
  wire [29:0] OptimizationBarrier_3_sum;
  wire [29:0] OptimizationBarrier_5_sum;
  wire [29:0] OptimizationBarrier_36_sum;
  wire [29:0] OptimizationBarrier_17_sum;
  wire [29:0] OptimizationBarrier_15_sum;
  wire [29:0] OptimizationBarrier_29_sum;
  wire [29:0] OptimizationBarrier_32_sum;
  wire [29:0] OptimizationBarrier_7_sum;
  wire [29:0] OptimizationBarrier_14_sum;
  wire [29:0] OptimizationBarrier_26_sum;
  wire [29:0] OptimizationBarrier_11_sum;
  wire [29:0] OptimizationBarrier_13_sum;
  wire  stopEn0;
  wire  OptimizationBarrier_34_metaAssert_wire;
  wire  OptimizationBarrier_20_metaAssert_wire;
  wire  OptimizationBarrier_6_metaAssert_wire;
  wire  OptimizationBarrier_22_metaAssert_wire;
  wire  OptimizationBarrier_14_metaAssert_wire;
  wire  OptimizationBarrier_36_metaAssert_wire;
  wire  OptimizationBarrier_37_metaAssert_wire;
  wire  OptimizationBarrier_16_metaAssert_wire;
  wire  OptimizationBarrier_35_metaAssert_wire;
  wire  OptimizationBarrier_metaAssert_wire;
  wire  OptimizationBarrier_24_metaAssert_wire;
  wire  OptimizationBarrier_32_metaAssert_wire;
  wire  pmp_metaAssert_wire;
  wire  OptimizationBarrier_33_metaAssert_wire;
  wire  OptimizationBarrier_25_metaAssert_wire;
  wire  OptimizationBarrier_4_metaAssert_wire;
  wire  OptimizationBarrier_30_metaAssert_wire;
  wire  OptimizationBarrier_23_metaAssert_wire;
  wire  OptimizationBarrier_7_metaAssert_wire;
  wire  OptimizationBarrier_10_metaAssert_wire;
  wire  OptimizationBarrier_15_metaAssert_wire;
  wire  OptimizationBarrier_8_metaAssert_wire;
  wire  OptimizationBarrier_28_metaAssert_wire;
  wire  OptimizationBarrier_3_metaAssert_wire;
  wire  OptimizationBarrier_18_metaAssert_wire;
  wire  OptimizationBarrier_2_metaAssert_wire;
  wire  OptimizationBarrier_31_metaAssert_wire;
  wire  OptimizationBarrier_26_metaAssert_wire;
  wire  OptimizationBarrier_11_metaAssert_wire;
  wire  OptimizationBarrier_19_metaAssert_wire;
  wire  OptimizationBarrier_9_metaAssert_wire;
  wire  OptimizationBarrier_1_metaAssert_wire;
  wire  OptimizationBarrier_5_metaAssert_wire;
  wire  OptimizationBarrier_12_metaAssert_wire;
  wire  OptimizationBarrier_38_metaAssert_wire;
  wire  OptimizationBarrier_17_metaAssert_wire;
  wire  OptimizationBarrier_27_metaAssert_wire;
  wire  OptimizationBarrier_29_metaAssert_wire;
  wire  OptimizationBarrier_13_metaAssert_wire;
  wire  OptimizationBarrier_21_metaAssert_wire;
  wire  TLB_or15;
  wire  TLB_or34;
  wire  TLB_or16;
  wire  TLB_or7;
  wire  TLB_or17;
  wire  TLB_or38;
  wire  TLB_or18;
  wire  TLB_or8;
  wire  TLB_or3;
  wire  TLB_or19;
  wire  TLB_or42;
  wire  TLB_or20;
  wire  TLB_or9;
  wire  TLB_or21;
  wire  TLB_or46;
  wire  TLB_or22;
  wire  TLB_or10;
  wire  TLB_or4;
  wire  TLB_or1;
  wire  TLB_or23;
  wire  TLB_or50;
  wire  TLB_or24;
  wire  TLB_or11;
  wire  TLB_or25;
  wire  TLB_or54;
  wire  TLB_or26;
  wire  TLB_or12;
  wire  TLB_or5;
  wire  TLB_or27;
  wire  TLB_or58;
  wire  TLB_or28;
  wire  TLB_or13;
  wire  TLB_or60;
  wire  TLB_or29;
  wire  TLB_or62;
  wire  TLB_or30;
  wire  TLB_or14;
  wire  TLB_or6;
  wire  TLB_or2;
  wire  TLB_or0;
  reg  TLB_metaAssert;
  reg [31:0] _RAND_103;
  OptimizationBarrier OptimizationBarrier ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_io_x_ppn),
    .io_x_u(OptimizationBarrier_io_x_u),
    .io_x_ae(OptimizationBarrier_io_x_ae),
    .io_x_sw(OptimizationBarrier_io_x_sw),
    .io_x_sx(OptimizationBarrier_io_x_sx),
    .io_x_sr(OptimizationBarrier_io_x_sr),
    .io_x_pw(OptimizationBarrier_io_x_pw),
    .io_x_px(OptimizationBarrier_io_x_px),
    .io_x_pr(OptimizationBarrier_io_x_pr),
    .io_x_ppp(OptimizationBarrier_io_x_ppp),
    .io_x_pal(OptimizationBarrier_io_x_pal),
    .io_x_paa(OptimizationBarrier_io_x_paa),
    .io_x_eff(OptimizationBarrier_io_x_eff),
    .io_x_c(OptimizationBarrier_io_x_c),
    .io_y_ppn(OptimizationBarrier_io_y_ppn),
    .io_y_u(OptimizationBarrier_io_y_u),
    .io_y_ae(OptimizationBarrier_io_y_ae),
    .io_y_sw(OptimizationBarrier_io_y_sw),
    .io_y_sx(OptimizationBarrier_io_y_sx),
    .io_y_sr(OptimizationBarrier_io_y_sr),
    .io_y_pw(OptimizationBarrier_io_y_pw),
    .io_y_px(OptimizationBarrier_io_y_px),
    .io_y_pr(OptimizationBarrier_io_y_pr),
    .io_y_ppp(OptimizationBarrier_io_y_ppp),
    .io_y_pal(OptimizationBarrier_io_y_pal),
    .io_y_paa(OptimizationBarrier_io_y_paa),
    .io_y_eff(OptimizationBarrier_io_y_eff),
    .io_y_c(OptimizationBarrier_io_y_c),
    .io_covSum(OptimizationBarrier_io_covSum),
    .metaAssert(OptimizationBarrier_metaAssert)
  );
  PMPChecker pmp ( // @[TLB.scala 190:19]
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_size(pmp_io_size),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x),
    .io_covSum(pmp_io_covSum),
    .metaAssert(pmp_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_1 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_1_io_x_ppn),
    .io_x_u(OptimizationBarrier_1_io_x_u),
    .io_x_ae(OptimizationBarrier_1_io_x_ae),
    .io_x_sw(OptimizationBarrier_1_io_x_sw),
    .io_x_sx(OptimizationBarrier_1_io_x_sx),
    .io_x_sr(OptimizationBarrier_1_io_x_sr),
    .io_x_pw(OptimizationBarrier_1_io_x_pw),
    .io_x_px(OptimizationBarrier_1_io_x_px),
    .io_x_pr(OptimizationBarrier_1_io_x_pr),
    .io_x_ppp(OptimizationBarrier_1_io_x_ppp),
    .io_x_pal(OptimizationBarrier_1_io_x_pal),
    .io_x_paa(OptimizationBarrier_1_io_x_paa),
    .io_x_eff(OptimizationBarrier_1_io_x_eff),
    .io_x_c(OptimizationBarrier_1_io_x_c),
    .io_y_ppn(OptimizationBarrier_1_io_y_ppn),
    .io_y_u(OptimizationBarrier_1_io_y_u),
    .io_y_ae(OptimizationBarrier_1_io_y_ae),
    .io_y_sw(OptimizationBarrier_1_io_y_sw),
    .io_y_sx(OptimizationBarrier_1_io_y_sx),
    .io_y_sr(OptimizationBarrier_1_io_y_sr),
    .io_y_pw(OptimizationBarrier_1_io_y_pw),
    .io_y_px(OptimizationBarrier_1_io_y_px),
    .io_y_pr(OptimizationBarrier_1_io_y_pr),
    .io_y_ppp(OptimizationBarrier_1_io_y_ppp),
    .io_y_pal(OptimizationBarrier_1_io_y_pal),
    .io_y_paa(OptimizationBarrier_1_io_y_paa),
    .io_y_eff(OptimizationBarrier_1_io_y_eff),
    .io_y_c(OptimizationBarrier_1_io_y_c),
    .io_covSum(OptimizationBarrier_1_io_covSum),
    .metaAssert(OptimizationBarrier_1_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_2 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_2_io_x_ppn),
    .io_x_u(OptimizationBarrier_2_io_x_u),
    .io_x_ae(OptimizationBarrier_2_io_x_ae),
    .io_x_sw(OptimizationBarrier_2_io_x_sw),
    .io_x_sx(OptimizationBarrier_2_io_x_sx),
    .io_x_sr(OptimizationBarrier_2_io_x_sr),
    .io_x_pw(OptimizationBarrier_2_io_x_pw),
    .io_x_px(OptimizationBarrier_2_io_x_px),
    .io_x_pr(OptimizationBarrier_2_io_x_pr),
    .io_x_ppp(OptimizationBarrier_2_io_x_ppp),
    .io_x_pal(OptimizationBarrier_2_io_x_pal),
    .io_x_paa(OptimizationBarrier_2_io_x_paa),
    .io_x_eff(OptimizationBarrier_2_io_x_eff),
    .io_x_c(OptimizationBarrier_2_io_x_c),
    .io_y_ppn(OptimizationBarrier_2_io_y_ppn),
    .io_y_u(OptimizationBarrier_2_io_y_u),
    .io_y_ae(OptimizationBarrier_2_io_y_ae),
    .io_y_sw(OptimizationBarrier_2_io_y_sw),
    .io_y_sx(OptimizationBarrier_2_io_y_sx),
    .io_y_sr(OptimizationBarrier_2_io_y_sr),
    .io_y_pw(OptimizationBarrier_2_io_y_pw),
    .io_y_px(OptimizationBarrier_2_io_y_px),
    .io_y_pr(OptimizationBarrier_2_io_y_pr),
    .io_y_ppp(OptimizationBarrier_2_io_y_ppp),
    .io_y_pal(OptimizationBarrier_2_io_y_pal),
    .io_y_paa(OptimizationBarrier_2_io_y_paa),
    .io_y_eff(OptimizationBarrier_2_io_y_eff),
    .io_y_c(OptimizationBarrier_2_io_y_c),
    .io_covSum(OptimizationBarrier_2_io_covSum),
    .metaAssert(OptimizationBarrier_2_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_3 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_3_io_x_ppn),
    .io_x_u(OptimizationBarrier_3_io_x_u),
    .io_x_ae(OptimizationBarrier_3_io_x_ae),
    .io_x_sw(OptimizationBarrier_3_io_x_sw),
    .io_x_sx(OptimizationBarrier_3_io_x_sx),
    .io_x_sr(OptimizationBarrier_3_io_x_sr),
    .io_x_pw(OptimizationBarrier_3_io_x_pw),
    .io_x_px(OptimizationBarrier_3_io_x_px),
    .io_x_pr(OptimizationBarrier_3_io_x_pr),
    .io_x_ppp(OptimizationBarrier_3_io_x_ppp),
    .io_x_pal(OptimizationBarrier_3_io_x_pal),
    .io_x_paa(OptimizationBarrier_3_io_x_paa),
    .io_x_eff(OptimizationBarrier_3_io_x_eff),
    .io_x_c(OptimizationBarrier_3_io_x_c),
    .io_y_ppn(OptimizationBarrier_3_io_y_ppn),
    .io_y_u(OptimizationBarrier_3_io_y_u),
    .io_y_ae(OptimizationBarrier_3_io_y_ae),
    .io_y_sw(OptimizationBarrier_3_io_y_sw),
    .io_y_sx(OptimizationBarrier_3_io_y_sx),
    .io_y_sr(OptimizationBarrier_3_io_y_sr),
    .io_y_pw(OptimizationBarrier_3_io_y_pw),
    .io_y_px(OptimizationBarrier_3_io_y_px),
    .io_y_pr(OptimizationBarrier_3_io_y_pr),
    .io_y_ppp(OptimizationBarrier_3_io_y_ppp),
    .io_y_pal(OptimizationBarrier_3_io_y_pal),
    .io_y_paa(OptimizationBarrier_3_io_y_paa),
    .io_y_eff(OptimizationBarrier_3_io_y_eff),
    .io_y_c(OptimizationBarrier_3_io_y_c),
    .io_covSum(OptimizationBarrier_3_io_covSum),
    .metaAssert(OptimizationBarrier_3_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_4 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_4_io_x_ppn),
    .io_x_u(OptimizationBarrier_4_io_x_u),
    .io_x_ae(OptimizationBarrier_4_io_x_ae),
    .io_x_sw(OptimizationBarrier_4_io_x_sw),
    .io_x_sx(OptimizationBarrier_4_io_x_sx),
    .io_x_sr(OptimizationBarrier_4_io_x_sr),
    .io_x_pw(OptimizationBarrier_4_io_x_pw),
    .io_x_px(OptimizationBarrier_4_io_x_px),
    .io_x_pr(OptimizationBarrier_4_io_x_pr),
    .io_x_ppp(OptimizationBarrier_4_io_x_ppp),
    .io_x_pal(OptimizationBarrier_4_io_x_pal),
    .io_x_paa(OptimizationBarrier_4_io_x_paa),
    .io_x_eff(OptimizationBarrier_4_io_x_eff),
    .io_x_c(OptimizationBarrier_4_io_x_c),
    .io_y_ppn(OptimizationBarrier_4_io_y_ppn),
    .io_y_u(OptimizationBarrier_4_io_y_u),
    .io_y_ae(OptimizationBarrier_4_io_y_ae),
    .io_y_sw(OptimizationBarrier_4_io_y_sw),
    .io_y_sx(OptimizationBarrier_4_io_y_sx),
    .io_y_sr(OptimizationBarrier_4_io_y_sr),
    .io_y_pw(OptimizationBarrier_4_io_y_pw),
    .io_y_px(OptimizationBarrier_4_io_y_px),
    .io_y_pr(OptimizationBarrier_4_io_y_pr),
    .io_y_ppp(OptimizationBarrier_4_io_y_ppp),
    .io_y_pal(OptimizationBarrier_4_io_y_pal),
    .io_y_paa(OptimizationBarrier_4_io_y_paa),
    .io_y_eff(OptimizationBarrier_4_io_y_eff),
    .io_y_c(OptimizationBarrier_4_io_y_c),
    .io_covSum(OptimizationBarrier_4_io_covSum),
    .metaAssert(OptimizationBarrier_4_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_5 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_5_io_x_ppn),
    .io_x_u(OptimizationBarrier_5_io_x_u),
    .io_x_ae(OptimizationBarrier_5_io_x_ae),
    .io_x_sw(OptimizationBarrier_5_io_x_sw),
    .io_x_sx(OptimizationBarrier_5_io_x_sx),
    .io_x_sr(OptimizationBarrier_5_io_x_sr),
    .io_x_pw(OptimizationBarrier_5_io_x_pw),
    .io_x_px(OptimizationBarrier_5_io_x_px),
    .io_x_pr(OptimizationBarrier_5_io_x_pr),
    .io_x_ppp(OptimizationBarrier_5_io_x_ppp),
    .io_x_pal(OptimizationBarrier_5_io_x_pal),
    .io_x_paa(OptimizationBarrier_5_io_x_paa),
    .io_x_eff(OptimizationBarrier_5_io_x_eff),
    .io_x_c(OptimizationBarrier_5_io_x_c),
    .io_y_ppn(OptimizationBarrier_5_io_y_ppn),
    .io_y_u(OptimizationBarrier_5_io_y_u),
    .io_y_ae(OptimizationBarrier_5_io_y_ae),
    .io_y_sw(OptimizationBarrier_5_io_y_sw),
    .io_y_sx(OptimizationBarrier_5_io_y_sx),
    .io_y_sr(OptimizationBarrier_5_io_y_sr),
    .io_y_pw(OptimizationBarrier_5_io_y_pw),
    .io_y_px(OptimizationBarrier_5_io_y_px),
    .io_y_pr(OptimizationBarrier_5_io_y_pr),
    .io_y_ppp(OptimizationBarrier_5_io_y_ppp),
    .io_y_pal(OptimizationBarrier_5_io_y_pal),
    .io_y_paa(OptimizationBarrier_5_io_y_paa),
    .io_y_eff(OptimizationBarrier_5_io_y_eff),
    .io_y_c(OptimizationBarrier_5_io_y_c),
    .io_covSum(OptimizationBarrier_5_io_covSum),
    .metaAssert(OptimizationBarrier_5_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_6 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_6_io_x_ppn),
    .io_x_u(OptimizationBarrier_6_io_x_u),
    .io_x_ae(OptimizationBarrier_6_io_x_ae),
    .io_x_sw(OptimizationBarrier_6_io_x_sw),
    .io_x_sx(OptimizationBarrier_6_io_x_sx),
    .io_x_sr(OptimizationBarrier_6_io_x_sr),
    .io_x_pw(OptimizationBarrier_6_io_x_pw),
    .io_x_px(OptimizationBarrier_6_io_x_px),
    .io_x_pr(OptimizationBarrier_6_io_x_pr),
    .io_x_ppp(OptimizationBarrier_6_io_x_ppp),
    .io_x_pal(OptimizationBarrier_6_io_x_pal),
    .io_x_paa(OptimizationBarrier_6_io_x_paa),
    .io_x_eff(OptimizationBarrier_6_io_x_eff),
    .io_x_c(OptimizationBarrier_6_io_x_c),
    .io_y_ppn(OptimizationBarrier_6_io_y_ppn),
    .io_y_u(OptimizationBarrier_6_io_y_u),
    .io_y_ae(OptimizationBarrier_6_io_y_ae),
    .io_y_sw(OptimizationBarrier_6_io_y_sw),
    .io_y_sx(OptimizationBarrier_6_io_y_sx),
    .io_y_sr(OptimizationBarrier_6_io_y_sr),
    .io_y_pw(OptimizationBarrier_6_io_y_pw),
    .io_y_px(OptimizationBarrier_6_io_y_px),
    .io_y_pr(OptimizationBarrier_6_io_y_pr),
    .io_y_ppp(OptimizationBarrier_6_io_y_ppp),
    .io_y_pal(OptimizationBarrier_6_io_y_pal),
    .io_y_paa(OptimizationBarrier_6_io_y_paa),
    .io_y_eff(OptimizationBarrier_6_io_y_eff),
    .io_y_c(OptimizationBarrier_6_io_y_c),
    .io_covSum(OptimizationBarrier_6_io_covSum),
    .metaAssert(OptimizationBarrier_6_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_7 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_7_io_x_ppn),
    .io_x_u(OptimizationBarrier_7_io_x_u),
    .io_x_ae(OptimizationBarrier_7_io_x_ae),
    .io_x_sw(OptimizationBarrier_7_io_x_sw),
    .io_x_sx(OptimizationBarrier_7_io_x_sx),
    .io_x_sr(OptimizationBarrier_7_io_x_sr),
    .io_x_pw(OptimizationBarrier_7_io_x_pw),
    .io_x_px(OptimizationBarrier_7_io_x_px),
    .io_x_pr(OptimizationBarrier_7_io_x_pr),
    .io_x_ppp(OptimizationBarrier_7_io_x_ppp),
    .io_x_pal(OptimizationBarrier_7_io_x_pal),
    .io_x_paa(OptimizationBarrier_7_io_x_paa),
    .io_x_eff(OptimizationBarrier_7_io_x_eff),
    .io_x_c(OptimizationBarrier_7_io_x_c),
    .io_y_ppn(OptimizationBarrier_7_io_y_ppn),
    .io_y_u(OptimizationBarrier_7_io_y_u),
    .io_y_ae(OptimizationBarrier_7_io_y_ae),
    .io_y_sw(OptimizationBarrier_7_io_y_sw),
    .io_y_sx(OptimizationBarrier_7_io_y_sx),
    .io_y_sr(OptimizationBarrier_7_io_y_sr),
    .io_y_pw(OptimizationBarrier_7_io_y_pw),
    .io_y_px(OptimizationBarrier_7_io_y_px),
    .io_y_pr(OptimizationBarrier_7_io_y_pr),
    .io_y_ppp(OptimizationBarrier_7_io_y_ppp),
    .io_y_pal(OptimizationBarrier_7_io_y_pal),
    .io_y_paa(OptimizationBarrier_7_io_y_paa),
    .io_y_eff(OptimizationBarrier_7_io_y_eff),
    .io_y_c(OptimizationBarrier_7_io_y_c),
    .io_covSum(OptimizationBarrier_7_io_covSum),
    .metaAssert(OptimizationBarrier_7_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_8 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_8_io_x_ppn),
    .io_x_u(OptimizationBarrier_8_io_x_u),
    .io_x_ae(OptimizationBarrier_8_io_x_ae),
    .io_x_sw(OptimizationBarrier_8_io_x_sw),
    .io_x_sx(OptimizationBarrier_8_io_x_sx),
    .io_x_sr(OptimizationBarrier_8_io_x_sr),
    .io_x_pw(OptimizationBarrier_8_io_x_pw),
    .io_x_px(OptimizationBarrier_8_io_x_px),
    .io_x_pr(OptimizationBarrier_8_io_x_pr),
    .io_x_ppp(OptimizationBarrier_8_io_x_ppp),
    .io_x_pal(OptimizationBarrier_8_io_x_pal),
    .io_x_paa(OptimizationBarrier_8_io_x_paa),
    .io_x_eff(OptimizationBarrier_8_io_x_eff),
    .io_x_c(OptimizationBarrier_8_io_x_c),
    .io_y_ppn(OptimizationBarrier_8_io_y_ppn),
    .io_y_u(OptimizationBarrier_8_io_y_u),
    .io_y_ae(OptimizationBarrier_8_io_y_ae),
    .io_y_sw(OptimizationBarrier_8_io_y_sw),
    .io_y_sx(OptimizationBarrier_8_io_y_sx),
    .io_y_sr(OptimizationBarrier_8_io_y_sr),
    .io_y_pw(OptimizationBarrier_8_io_y_pw),
    .io_y_px(OptimizationBarrier_8_io_y_px),
    .io_y_pr(OptimizationBarrier_8_io_y_pr),
    .io_y_ppp(OptimizationBarrier_8_io_y_ppp),
    .io_y_pal(OptimizationBarrier_8_io_y_pal),
    .io_y_paa(OptimizationBarrier_8_io_y_paa),
    .io_y_eff(OptimizationBarrier_8_io_y_eff),
    .io_y_c(OptimizationBarrier_8_io_y_c),
    .io_covSum(OptimizationBarrier_8_io_covSum),
    .metaAssert(OptimizationBarrier_8_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_9 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_9_io_x_ppn),
    .io_x_u(OptimizationBarrier_9_io_x_u),
    .io_x_ae(OptimizationBarrier_9_io_x_ae),
    .io_x_sw(OptimizationBarrier_9_io_x_sw),
    .io_x_sx(OptimizationBarrier_9_io_x_sx),
    .io_x_sr(OptimizationBarrier_9_io_x_sr),
    .io_x_pw(OptimizationBarrier_9_io_x_pw),
    .io_x_px(OptimizationBarrier_9_io_x_px),
    .io_x_pr(OptimizationBarrier_9_io_x_pr),
    .io_x_ppp(OptimizationBarrier_9_io_x_ppp),
    .io_x_pal(OptimizationBarrier_9_io_x_pal),
    .io_x_paa(OptimizationBarrier_9_io_x_paa),
    .io_x_eff(OptimizationBarrier_9_io_x_eff),
    .io_x_c(OptimizationBarrier_9_io_x_c),
    .io_y_ppn(OptimizationBarrier_9_io_y_ppn),
    .io_y_u(OptimizationBarrier_9_io_y_u),
    .io_y_ae(OptimizationBarrier_9_io_y_ae),
    .io_y_sw(OptimizationBarrier_9_io_y_sw),
    .io_y_sx(OptimizationBarrier_9_io_y_sx),
    .io_y_sr(OptimizationBarrier_9_io_y_sr),
    .io_y_pw(OptimizationBarrier_9_io_y_pw),
    .io_y_px(OptimizationBarrier_9_io_y_px),
    .io_y_pr(OptimizationBarrier_9_io_y_pr),
    .io_y_ppp(OptimizationBarrier_9_io_y_ppp),
    .io_y_pal(OptimizationBarrier_9_io_y_pal),
    .io_y_paa(OptimizationBarrier_9_io_y_paa),
    .io_y_eff(OptimizationBarrier_9_io_y_eff),
    .io_y_c(OptimizationBarrier_9_io_y_c),
    .io_covSum(OptimizationBarrier_9_io_covSum),
    .metaAssert(OptimizationBarrier_9_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_10 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_10_io_x_ppn),
    .io_x_u(OptimizationBarrier_10_io_x_u),
    .io_x_ae(OptimizationBarrier_10_io_x_ae),
    .io_x_sw(OptimizationBarrier_10_io_x_sw),
    .io_x_sx(OptimizationBarrier_10_io_x_sx),
    .io_x_sr(OptimizationBarrier_10_io_x_sr),
    .io_x_pw(OptimizationBarrier_10_io_x_pw),
    .io_x_px(OptimizationBarrier_10_io_x_px),
    .io_x_pr(OptimizationBarrier_10_io_x_pr),
    .io_x_ppp(OptimizationBarrier_10_io_x_ppp),
    .io_x_pal(OptimizationBarrier_10_io_x_pal),
    .io_x_paa(OptimizationBarrier_10_io_x_paa),
    .io_x_eff(OptimizationBarrier_10_io_x_eff),
    .io_x_c(OptimizationBarrier_10_io_x_c),
    .io_y_ppn(OptimizationBarrier_10_io_y_ppn),
    .io_y_u(OptimizationBarrier_10_io_y_u),
    .io_y_ae(OptimizationBarrier_10_io_y_ae),
    .io_y_sw(OptimizationBarrier_10_io_y_sw),
    .io_y_sx(OptimizationBarrier_10_io_y_sx),
    .io_y_sr(OptimizationBarrier_10_io_y_sr),
    .io_y_pw(OptimizationBarrier_10_io_y_pw),
    .io_y_px(OptimizationBarrier_10_io_y_px),
    .io_y_pr(OptimizationBarrier_10_io_y_pr),
    .io_y_ppp(OptimizationBarrier_10_io_y_ppp),
    .io_y_pal(OptimizationBarrier_10_io_y_pal),
    .io_y_paa(OptimizationBarrier_10_io_y_paa),
    .io_y_eff(OptimizationBarrier_10_io_y_eff),
    .io_y_c(OptimizationBarrier_10_io_y_c),
    .io_covSum(OptimizationBarrier_10_io_covSum),
    .metaAssert(OptimizationBarrier_10_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_11 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_11_io_x_ppn),
    .io_x_u(OptimizationBarrier_11_io_x_u),
    .io_x_ae(OptimizationBarrier_11_io_x_ae),
    .io_x_sw(OptimizationBarrier_11_io_x_sw),
    .io_x_sx(OptimizationBarrier_11_io_x_sx),
    .io_x_sr(OptimizationBarrier_11_io_x_sr),
    .io_x_pw(OptimizationBarrier_11_io_x_pw),
    .io_x_px(OptimizationBarrier_11_io_x_px),
    .io_x_pr(OptimizationBarrier_11_io_x_pr),
    .io_x_ppp(OptimizationBarrier_11_io_x_ppp),
    .io_x_pal(OptimizationBarrier_11_io_x_pal),
    .io_x_paa(OptimizationBarrier_11_io_x_paa),
    .io_x_eff(OptimizationBarrier_11_io_x_eff),
    .io_x_c(OptimizationBarrier_11_io_x_c),
    .io_y_ppn(OptimizationBarrier_11_io_y_ppn),
    .io_y_u(OptimizationBarrier_11_io_y_u),
    .io_y_ae(OptimizationBarrier_11_io_y_ae),
    .io_y_sw(OptimizationBarrier_11_io_y_sw),
    .io_y_sx(OptimizationBarrier_11_io_y_sx),
    .io_y_sr(OptimizationBarrier_11_io_y_sr),
    .io_y_pw(OptimizationBarrier_11_io_y_pw),
    .io_y_px(OptimizationBarrier_11_io_y_px),
    .io_y_pr(OptimizationBarrier_11_io_y_pr),
    .io_y_ppp(OptimizationBarrier_11_io_y_ppp),
    .io_y_pal(OptimizationBarrier_11_io_y_pal),
    .io_y_paa(OptimizationBarrier_11_io_y_paa),
    .io_y_eff(OptimizationBarrier_11_io_y_eff),
    .io_y_c(OptimizationBarrier_11_io_y_c),
    .io_covSum(OptimizationBarrier_11_io_covSum),
    .metaAssert(OptimizationBarrier_11_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_12 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_12_io_x_ppn),
    .io_x_u(OptimizationBarrier_12_io_x_u),
    .io_x_ae(OptimizationBarrier_12_io_x_ae),
    .io_x_sw(OptimizationBarrier_12_io_x_sw),
    .io_x_sx(OptimizationBarrier_12_io_x_sx),
    .io_x_sr(OptimizationBarrier_12_io_x_sr),
    .io_x_pw(OptimizationBarrier_12_io_x_pw),
    .io_x_px(OptimizationBarrier_12_io_x_px),
    .io_x_pr(OptimizationBarrier_12_io_x_pr),
    .io_x_ppp(OptimizationBarrier_12_io_x_ppp),
    .io_x_pal(OptimizationBarrier_12_io_x_pal),
    .io_x_paa(OptimizationBarrier_12_io_x_paa),
    .io_x_eff(OptimizationBarrier_12_io_x_eff),
    .io_x_c(OptimizationBarrier_12_io_x_c),
    .io_y_ppn(OptimizationBarrier_12_io_y_ppn),
    .io_y_u(OptimizationBarrier_12_io_y_u),
    .io_y_ae(OptimizationBarrier_12_io_y_ae),
    .io_y_sw(OptimizationBarrier_12_io_y_sw),
    .io_y_sx(OptimizationBarrier_12_io_y_sx),
    .io_y_sr(OptimizationBarrier_12_io_y_sr),
    .io_y_pw(OptimizationBarrier_12_io_y_pw),
    .io_y_px(OptimizationBarrier_12_io_y_px),
    .io_y_pr(OptimizationBarrier_12_io_y_pr),
    .io_y_ppp(OptimizationBarrier_12_io_y_ppp),
    .io_y_pal(OptimizationBarrier_12_io_y_pal),
    .io_y_paa(OptimizationBarrier_12_io_y_paa),
    .io_y_eff(OptimizationBarrier_12_io_y_eff),
    .io_y_c(OptimizationBarrier_12_io_y_c),
    .io_covSum(OptimizationBarrier_12_io_covSum),
    .metaAssert(OptimizationBarrier_12_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_13 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_13_io_x_ppn),
    .io_x_u(OptimizationBarrier_13_io_x_u),
    .io_x_ae(OptimizationBarrier_13_io_x_ae),
    .io_x_sw(OptimizationBarrier_13_io_x_sw),
    .io_x_sx(OptimizationBarrier_13_io_x_sx),
    .io_x_sr(OptimizationBarrier_13_io_x_sr),
    .io_x_pw(OptimizationBarrier_13_io_x_pw),
    .io_x_px(OptimizationBarrier_13_io_x_px),
    .io_x_pr(OptimizationBarrier_13_io_x_pr),
    .io_x_ppp(OptimizationBarrier_13_io_x_ppp),
    .io_x_pal(OptimizationBarrier_13_io_x_pal),
    .io_x_paa(OptimizationBarrier_13_io_x_paa),
    .io_x_eff(OptimizationBarrier_13_io_x_eff),
    .io_x_c(OptimizationBarrier_13_io_x_c),
    .io_y_ppn(OptimizationBarrier_13_io_y_ppn),
    .io_y_u(OptimizationBarrier_13_io_y_u),
    .io_y_ae(OptimizationBarrier_13_io_y_ae),
    .io_y_sw(OptimizationBarrier_13_io_y_sw),
    .io_y_sx(OptimizationBarrier_13_io_y_sx),
    .io_y_sr(OptimizationBarrier_13_io_y_sr),
    .io_y_pw(OptimizationBarrier_13_io_y_pw),
    .io_y_px(OptimizationBarrier_13_io_y_px),
    .io_y_pr(OptimizationBarrier_13_io_y_pr),
    .io_y_ppp(OptimizationBarrier_13_io_y_ppp),
    .io_y_pal(OptimizationBarrier_13_io_y_pal),
    .io_y_paa(OptimizationBarrier_13_io_y_paa),
    .io_y_eff(OptimizationBarrier_13_io_y_eff),
    .io_y_c(OptimizationBarrier_13_io_y_c),
    .io_covSum(OptimizationBarrier_13_io_covSum),
    .metaAssert(OptimizationBarrier_13_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_14 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_14_io_x_ppn),
    .io_x_u(OptimizationBarrier_14_io_x_u),
    .io_x_ae(OptimizationBarrier_14_io_x_ae),
    .io_x_sw(OptimizationBarrier_14_io_x_sw),
    .io_x_sx(OptimizationBarrier_14_io_x_sx),
    .io_x_sr(OptimizationBarrier_14_io_x_sr),
    .io_x_pw(OptimizationBarrier_14_io_x_pw),
    .io_x_px(OptimizationBarrier_14_io_x_px),
    .io_x_pr(OptimizationBarrier_14_io_x_pr),
    .io_x_ppp(OptimizationBarrier_14_io_x_ppp),
    .io_x_pal(OptimizationBarrier_14_io_x_pal),
    .io_x_paa(OptimizationBarrier_14_io_x_paa),
    .io_x_eff(OptimizationBarrier_14_io_x_eff),
    .io_x_c(OptimizationBarrier_14_io_x_c),
    .io_y_ppn(OptimizationBarrier_14_io_y_ppn),
    .io_y_u(OptimizationBarrier_14_io_y_u),
    .io_y_ae(OptimizationBarrier_14_io_y_ae),
    .io_y_sw(OptimizationBarrier_14_io_y_sw),
    .io_y_sx(OptimizationBarrier_14_io_y_sx),
    .io_y_sr(OptimizationBarrier_14_io_y_sr),
    .io_y_pw(OptimizationBarrier_14_io_y_pw),
    .io_y_px(OptimizationBarrier_14_io_y_px),
    .io_y_pr(OptimizationBarrier_14_io_y_pr),
    .io_y_ppp(OptimizationBarrier_14_io_y_ppp),
    .io_y_pal(OptimizationBarrier_14_io_y_pal),
    .io_y_paa(OptimizationBarrier_14_io_y_paa),
    .io_y_eff(OptimizationBarrier_14_io_y_eff),
    .io_y_c(OptimizationBarrier_14_io_y_c),
    .io_covSum(OptimizationBarrier_14_io_covSum),
    .metaAssert(OptimizationBarrier_14_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_15 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_15_io_x_ppn),
    .io_x_u(OptimizationBarrier_15_io_x_u),
    .io_x_ae(OptimizationBarrier_15_io_x_ae),
    .io_x_sw(OptimizationBarrier_15_io_x_sw),
    .io_x_sx(OptimizationBarrier_15_io_x_sx),
    .io_x_sr(OptimizationBarrier_15_io_x_sr),
    .io_x_pw(OptimizationBarrier_15_io_x_pw),
    .io_x_px(OptimizationBarrier_15_io_x_px),
    .io_x_pr(OptimizationBarrier_15_io_x_pr),
    .io_x_ppp(OptimizationBarrier_15_io_x_ppp),
    .io_x_pal(OptimizationBarrier_15_io_x_pal),
    .io_x_paa(OptimizationBarrier_15_io_x_paa),
    .io_x_eff(OptimizationBarrier_15_io_x_eff),
    .io_x_c(OptimizationBarrier_15_io_x_c),
    .io_y_ppn(OptimizationBarrier_15_io_y_ppn),
    .io_y_u(OptimizationBarrier_15_io_y_u),
    .io_y_ae(OptimizationBarrier_15_io_y_ae),
    .io_y_sw(OptimizationBarrier_15_io_y_sw),
    .io_y_sx(OptimizationBarrier_15_io_y_sx),
    .io_y_sr(OptimizationBarrier_15_io_y_sr),
    .io_y_pw(OptimizationBarrier_15_io_y_pw),
    .io_y_px(OptimizationBarrier_15_io_y_px),
    .io_y_pr(OptimizationBarrier_15_io_y_pr),
    .io_y_ppp(OptimizationBarrier_15_io_y_ppp),
    .io_y_pal(OptimizationBarrier_15_io_y_pal),
    .io_y_paa(OptimizationBarrier_15_io_y_paa),
    .io_y_eff(OptimizationBarrier_15_io_y_eff),
    .io_y_c(OptimizationBarrier_15_io_y_c),
    .io_covSum(OptimizationBarrier_15_io_covSum),
    .metaAssert(OptimizationBarrier_15_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_16 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_16_io_x_ppn),
    .io_x_u(OptimizationBarrier_16_io_x_u),
    .io_x_ae(OptimizationBarrier_16_io_x_ae),
    .io_x_sw(OptimizationBarrier_16_io_x_sw),
    .io_x_sx(OptimizationBarrier_16_io_x_sx),
    .io_x_sr(OptimizationBarrier_16_io_x_sr),
    .io_x_pw(OptimizationBarrier_16_io_x_pw),
    .io_x_px(OptimizationBarrier_16_io_x_px),
    .io_x_pr(OptimizationBarrier_16_io_x_pr),
    .io_x_ppp(OptimizationBarrier_16_io_x_ppp),
    .io_x_pal(OptimizationBarrier_16_io_x_pal),
    .io_x_paa(OptimizationBarrier_16_io_x_paa),
    .io_x_eff(OptimizationBarrier_16_io_x_eff),
    .io_x_c(OptimizationBarrier_16_io_x_c),
    .io_y_ppn(OptimizationBarrier_16_io_y_ppn),
    .io_y_u(OptimizationBarrier_16_io_y_u),
    .io_y_ae(OptimizationBarrier_16_io_y_ae),
    .io_y_sw(OptimizationBarrier_16_io_y_sw),
    .io_y_sx(OptimizationBarrier_16_io_y_sx),
    .io_y_sr(OptimizationBarrier_16_io_y_sr),
    .io_y_pw(OptimizationBarrier_16_io_y_pw),
    .io_y_px(OptimizationBarrier_16_io_y_px),
    .io_y_pr(OptimizationBarrier_16_io_y_pr),
    .io_y_ppp(OptimizationBarrier_16_io_y_ppp),
    .io_y_pal(OptimizationBarrier_16_io_y_pal),
    .io_y_paa(OptimizationBarrier_16_io_y_paa),
    .io_y_eff(OptimizationBarrier_16_io_y_eff),
    .io_y_c(OptimizationBarrier_16_io_y_c),
    .io_covSum(OptimizationBarrier_16_io_covSum),
    .metaAssert(OptimizationBarrier_16_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_17 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_17_io_x_ppn),
    .io_x_u(OptimizationBarrier_17_io_x_u),
    .io_x_ae(OptimizationBarrier_17_io_x_ae),
    .io_x_sw(OptimizationBarrier_17_io_x_sw),
    .io_x_sx(OptimizationBarrier_17_io_x_sx),
    .io_x_sr(OptimizationBarrier_17_io_x_sr),
    .io_x_pw(OptimizationBarrier_17_io_x_pw),
    .io_x_px(OptimizationBarrier_17_io_x_px),
    .io_x_pr(OptimizationBarrier_17_io_x_pr),
    .io_x_ppp(OptimizationBarrier_17_io_x_ppp),
    .io_x_pal(OptimizationBarrier_17_io_x_pal),
    .io_x_paa(OptimizationBarrier_17_io_x_paa),
    .io_x_eff(OptimizationBarrier_17_io_x_eff),
    .io_x_c(OptimizationBarrier_17_io_x_c),
    .io_y_ppn(OptimizationBarrier_17_io_y_ppn),
    .io_y_u(OptimizationBarrier_17_io_y_u),
    .io_y_ae(OptimizationBarrier_17_io_y_ae),
    .io_y_sw(OptimizationBarrier_17_io_y_sw),
    .io_y_sx(OptimizationBarrier_17_io_y_sx),
    .io_y_sr(OptimizationBarrier_17_io_y_sr),
    .io_y_pw(OptimizationBarrier_17_io_y_pw),
    .io_y_px(OptimizationBarrier_17_io_y_px),
    .io_y_pr(OptimizationBarrier_17_io_y_pr),
    .io_y_ppp(OptimizationBarrier_17_io_y_ppp),
    .io_y_pal(OptimizationBarrier_17_io_y_pal),
    .io_y_paa(OptimizationBarrier_17_io_y_paa),
    .io_y_eff(OptimizationBarrier_17_io_y_eff),
    .io_y_c(OptimizationBarrier_17_io_y_c),
    .io_covSum(OptimizationBarrier_17_io_covSum),
    .metaAssert(OptimizationBarrier_17_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_18 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_18_io_x_ppn),
    .io_x_u(OptimizationBarrier_18_io_x_u),
    .io_x_ae(OptimizationBarrier_18_io_x_ae),
    .io_x_sw(OptimizationBarrier_18_io_x_sw),
    .io_x_sx(OptimizationBarrier_18_io_x_sx),
    .io_x_sr(OptimizationBarrier_18_io_x_sr),
    .io_x_pw(OptimizationBarrier_18_io_x_pw),
    .io_x_px(OptimizationBarrier_18_io_x_px),
    .io_x_pr(OptimizationBarrier_18_io_x_pr),
    .io_x_ppp(OptimizationBarrier_18_io_x_ppp),
    .io_x_pal(OptimizationBarrier_18_io_x_pal),
    .io_x_paa(OptimizationBarrier_18_io_x_paa),
    .io_x_eff(OptimizationBarrier_18_io_x_eff),
    .io_x_c(OptimizationBarrier_18_io_x_c),
    .io_y_ppn(OptimizationBarrier_18_io_y_ppn),
    .io_y_u(OptimizationBarrier_18_io_y_u),
    .io_y_ae(OptimizationBarrier_18_io_y_ae),
    .io_y_sw(OptimizationBarrier_18_io_y_sw),
    .io_y_sx(OptimizationBarrier_18_io_y_sx),
    .io_y_sr(OptimizationBarrier_18_io_y_sr),
    .io_y_pw(OptimizationBarrier_18_io_y_pw),
    .io_y_px(OptimizationBarrier_18_io_y_px),
    .io_y_pr(OptimizationBarrier_18_io_y_pr),
    .io_y_ppp(OptimizationBarrier_18_io_y_ppp),
    .io_y_pal(OptimizationBarrier_18_io_y_pal),
    .io_y_paa(OptimizationBarrier_18_io_y_paa),
    .io_y_eff(OptimizationBarrier_18_io_y_eff),
    .io_y_c(OptimizationBarrier_18_io_y_c),
    .io_covSum(OptimizationBarrier_18_io_covSum),
    .metaAssert(OptimizationBarrier_18_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_19 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_19_io_x_ppn),
    .io_x_u(OptimizationBarrier_19_io_x_u),
    .io_x_ae(OptimizationBarrier_19_io_x_ae),
    .io_x_sw(OptimizationBarrier_19_io_x_sw),
    .io_x_sx(OptimizationBarrier_19_io_x_sx),
    .io_x_sr(OptimizationBarrier_19_io_x_sr),
    .io_x_pw(OptimizationBarrier_19_io_x_pw),
    .io_x_px(OptimizationBarrier_19_io_x_px),
    .io_x_pr(OptimizationBarrier_19_io_x_pr),
    .io_x_ppp(OptimizationBarrier_19_io_x_ppp),
    .io_x_pal(OptimizationBarrier_19_io_x_pal),
    .io_x_paa(OptimizationBarrier_19_io_x_paa),
    .io_x_eff(OptimizationBarrier_19_io_x_eff),
    .io_x_c(OptimizationBarrier_19_io_x_c),
    .io_y_ppn(OptimizationBarrier_19_io_y_ppn),
    .io_y_u(OptimizationBarrier_19_io_y_u),
    .io_y_ae(OptimizationBarrier_19_io_y_ae),
    .io_y_sw(OptimizationBarrier_19_io_y_sw),
    .io_y_sx(OptimizationBarrier_19_io_y_sx),
    .io_y_sr(OptimizationBarrier_19_io_y_sr),
    .io_y_pw(OptimizationBarrier_19_io_y_pw),
    .io_y_px(OptimizationBarrier_19_io_y_px),
    .io_y_pr(OptimizationBarrier_19_io_y_pr),
    .io_y_ppp(OptimizationBarrier_19_io_y_ppp),
    .io_y_pal(OptimizationBarrier_19_io_y_pal),
    .io_y_paa(OptimizationBarrier_19_io_y_paa),
    .io_y_eff(OptimizationBarrier_19_io_y_eff),
    .io_y_c(OptimizationBarrier_19_io_y_c),
    .io_covSum(OptimizationBarrier_19_io_covSum),
    .metaAssert(OptimizationBarrier_19_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_20 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_20_io_x_ppn),
    .io_x_u(OptimizationBarrier_20_io_x_u),
    .io_x_ae(OptimizationBarrier_20_io_x_ae),
    .io_x_sw(OptimizationBarrier_20_io_x_sw),
    .io_x_sx(OptimizationBarrier_20_io_x_sx),
    .io_x_sr(OptimizationBarrier_20_io_x_sr),
    .io_x_pw(OptimizationBarrier_20_io_x_pw),
    .io_x_px(OptimizationBarrier_20_io_x_px),
    .io_x_pr(OptimizationBarrier_20_io_x_pr),
    .io_x_ppp(OptimizationBarrier_20_io_x_ppp),
    .io_x_pal(OptimizationBarrier_20_io_x_pal),
    .io_x_paa(OptimizationBarrier_20_io_x_paa),
    .io_x_eff(OptimizationBarrier_20_io_x_eff),
    .io_x_c(OptimizationBarrier_20_io_x_c),
    .io_y_ppn(OptimizationBarrier_20_io_y_ppn),
    .io_y_u(OptimizationBarrier_20_io_y_u),
    .io_y_ae(OptimizationBarrier_20_io_y_ae),
    .io_y_sw(OptimizationBarrier_20_io_y_sw),
    .io_y_sx(OptimizationBarrier_20_io_y_sx),
    .io_y_sr(OptimizationBarrier_20_io_y_sr),
    .io_y_pw(OptimizationBarrier_20_io_y_pw),
    .io_y_px(OptimizationBarrier_20_io_y_px),
    .io_y_pr(OptimizationBarrier_20_io_y_pr),
    .io_y_ppp(OptimizationBarrier_20_io_y_ppp),
    .io_y_pal(OptimizationBarrier_20_io_y_pal),
    .io_y_paa(OptimizationBarrier_20_io_y_paa),
    .io_y_eff(OptimizationBarrier_20_io_y_eff),
    .io_y_c(OptimizationBarrier_20_io_y_c),
    .io_covSum(OptimizationBarrier_20_io_covSum),
    .metaAssert(OptimizationBarrier_20_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_21 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_21_io_x_ppn),
    .io_x_u(OptimizationBarrier_21_io_x_u),
    .io_x_ae(OptimizationBarrier_21_io_x_ae),
    .io_x_sw(OptimizationBarrier_21_io_x_sw),
    .io_x_sx(OptimizationBarrier_21_io_x_sx),
    .io_x_sr(OptimizationBarrier_21_io_x_sr),
    .io_x_pw(OptimizationBarrier_21_io_x_pw),
    .io_x_px(OptimizationBarrier_21_io_x_px),
    .io_x_pr(OptimizationBarrier_21_io_x_pr),
    .io_x_ppp(OptimizationBarrier_21_io_x_ppp),
    .io_x_pal(OptimizationBarrier_21_io_x_pal),
    .io_x_paa(OptimizationBarrier_21_io_x_paa),
    .io_x_eff(OptimizationBarrier_21_io_x_eff),
    .io_x_c(OptimizationBarrier_21_io_x_c),
    .io_y_ppn(OptimizationBarrier_21_io_y_ppn),
    .io_y_u(OptimizationBarrier_21_io_y_u),
    .io_y_ae(OptimizationBarrier_21_io_y_ae),
    .io_y_sw(OptimizationBarrier_21_io_y_sw),
    .io_y_sx(OptimizationBarrier_21_io_y_sx),
    .io_y_sr(OptimizationBarrier_21_io_y_sr),
    .io_y_pw(OptimizationBarrier_21_io_y_pw),
    .io_y_px(OptimizationBarrier_21_io_y_px),
    .io_y_pr(OptimizationBarrier_21_io_y_pr),
    .io_y_ppp(OptimizationBarrier_21_io_y_ppp),
    .io_y_pal(OptimizationBarrier_21_io_y_pal),
    .io_y_paa(OptimizationBarrier_21_io_y_paa),
    .io_y_eff(OptimizationBarrier_21_io_y_eff),
    .io_y_c(OptimizationBarrier_21_io_y_c),
    .io_covSum(OptimizationBarrier_21_io_covSum),
    .metaAssert(OptimizationBarrier_21_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_22 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_22_io_x_ppn),
    .io_x_u(OptimizationBarrier_22_io_x_u),
    .io_x_ae(OptimizationBarrier_22_io_x_ae),
    .io_x_sw(OptimizationBarrier_22_io_x_sw),
    .io_x_sx(OptimizationBarrier_22_io_x_sx),
    .io_x_sr(OptimizationBarrier_22_io_x_sr),
    .io_x_pw(OptimizationBarrier_22_io_x_pw),
    .io_x_px(OptimizationBarrier_22_io_x_px),
    .io_x_pr(OptimizationBarrier_22_io_x_pr),
    .io_x_ppp(OptimizationBarrier_22_io_x_ppp),
    .io_x_pal(OptimizationBarrier_22_io_x_pal),
    .io_x_paa(OptimizationBarrier_22_io_x_paa),
    .io_x_eff(OptimizationBarrier_22_io_x_eff),
    .io_x_c(OptimizationBarrier_22_io_x_c),
    .io_y_ppn(OptimizationBarrier_22_io_y_ppn),
    .io_y_u(OptimizationBarrier_22_io_y_u),
    .io_y_ae(OptimizationBarrier_22_io_y_ae),
    .io_y_sw(OptimizationBarrier_22_io_y_sw),
    .io_y_sx(OptimizationBarrier_22_io_y_sx),
    .io_y_sr(OptimizationBarrier_22_io_y_sr),
    .io_y_pw(OptimizationBarrier_22_io_y_pw),
    .io_y_px(OptimizationBarrier_22_io_y_px),
    .io_y_pr(OptimizationBarrier_22_io_y_pr),
    .io_y_ppp(OptimizationBarrier_22_io_y_ppp),
    .io_y_pal(OptimizationBarrier_22_io_y_pal),
    .io_y_paa(OptimizationBarrier_22_io_y_paa),
    .io_y_eff(OptimizationBarrier_22_io_y_eff),
    .io_y_c(OptimizationBarrier_22_io_y_c),
    .io_covSum(OptimizationBarrier_22_io_covSum),
    .metaAssert(OptimizationBarrier_22_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_23 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_23_io_x_ppn),
    .io_x_u(OptimizationBarrier_23_io_x_u),
    .io_x_ae(OptimizationBarrier_23_io_x_ae),
    .io_x_sw(OptimizationBarrier_23_io_x_sw),
    .io_x_sx(OptimizationBarrier_23_io_x_sx),
    .io_x_sr(OptimizationBarrier_23_io_x_sr),
    .io_x_pw(OptimizationBarrier_23_io_x_pw),
    .io_x_px(OptimizationBarrier_23_io_x_px),
    .io_x_pr(OptimizationBarrier_23_io_x_pr),
    .io_x_ppp(OptimizationBarrier_23_io_x_ppp),
    .io_x_pal(OptimizationBarrier_23_io_x_pal),
    .io_x_paa(OptimizationBarrier_23_io_x_paa),
    .io_x_eff(OptimizationBarrier_23_io_x_eff),
    .io_x_c(OptimizationBarrier_23_io_x_c),
    .io_y_ppn(OptimizationBarrier_23_io_y_ppn),
    .io_y_u(OptimizationBarrier_23_io_y_u),
    .io_y_ae(OptimizationBarrier_23_io_y_ae),
    .io_y_sw(OptimizationBarrier_23_io_y_sw),
    .io_y_sx(OptimizationBarrier_23_io_y_sx),
    .io_y_sr(OptimizationBarrier_23_io_y_sr),
    .io_y_pw(OptimizationBarrier_23_io_y_pw),
    .io_y_px(OptimizationBarrier_23_io_y_px),
    .io_y_pr(OptimizationBarrier_23_io_y_pr),
    .io_y_ppp(OptimizationBarrier_23_io_y_ppp),
    .io_y_pal(OptimizationBarrier_23_io_y_pal),
    .io_y_paa(OptimizationBarrier_23_io_y_paa),
    .io_y_eff(OptimizationBarrier_23_io_y_eff),
    .io_y_c(OptimizationBarrier_23_io_y_c),
    .io_covSum(OptimizationBarrier_23_io_covSum),
    .metaAssert(OptimizationBarrier_23_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_24 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_24_io_x_ppn),
    .io_x_u(OptimizationBarrier_24_io_x_u),
    .io_x_ae(OptimizationBarrier_24_io_x_ae),
    .io_x_sw(OptimizationBarrier_24_io_x_sw),
    .io_x_sx(OptimizationBarrier_24_io_x_sx),
    .io_x_sr(OptimizationBarrier_24_io_x_sr),
    .io_x_pw(OptimizationBarrier_24_io_x_pw),
    .io_x_px(OptimizationBarrier_24_io_x_px),
    .io_x_pr(OptimizationBarrier_24_io_x_pr),
    .io_x_ppp(OptimizationBarrier_24_io_x_ppp),
    .io_x_pal(OptimizationBarrier_24_io_x_pal),
    .io_x_paa(OptimizationBarrier_24_io_x_paa),
    .io_x_eff(OptimizationBarrier_24_io_x_eff),
    .io_x_c(OptimizationBarrier_24_io_x_c),
    .io_y_ppn(OptimizationBarrier_24_io_y_ppn),
    .io_y_u(OptimizationBarrier_24_io_y_u),
    .io_y_ae(OptimizationBarrier_24_io_y_ae),
    .io_y_sw(OptimizationBarrier_24_io_y_sw),
    .io_y_sx(OptimizationBarrier_24_io_y_sx),
    .io_y_sr(OptimizationBarrier_24_io_y_sr),
    .io_y_pw(OptimizationBarrier_24_io_y_pw),
    .io_y_px(OptimizationBarrier_24_io_y_px),
    .io_y_pr(OptimizationBarrier_24_io_y_pr),
    .io_y_ppp(OptimizationBarrier_24_io_y_ppp),
    .io_y_pal(OptimizationBarrier_24_io_y_pal),
    .io_y_paa(OptimizationBarrier_24_io_y_paa),
    .io_y_eff(OptimizationBarrier_24_io_y_eff),
    .io_y_c(OptimizationBarrier_24_io_y_c),
    .io_covSum(OptimizationBarrier_24_io_covSum),
    .metaAssert(OptimizationBarrier_24_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_25 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_25_io_x_ppn),
    .io_x_u(OptimizationBarrier_25_io_x_u),
    .io_x_ae(OptimizationBarrier_25_io_x_ae),
    .io_x_sw(OptimizationBarrier_25_io_x_sw),
    .io_x_sx(OptimizationBarrier_25_io_x_sx),
    .io_x_sr(OptimizationBarrier_25_io_x_sr),
    .io_x_pw(OptimizationBarrier_25_io_x_pw),
    .io_x_px(OptimizationBarrier_25_io_x_px),
    .io_x_pr(OptimizationBarrier_25_io_x_pr),
    .io_x_ppp(OptimizationBarrier_25_io_x_ppp),
    .io_x_pal(OptimizationBarrier_25_io_x_pal),
    .io_x_paa(OptimizationBarrier_25_io_x_paa),
    .io_x_eff(OptimizationBarrier_25_io_x_eff),
    .io_x_c(OptimizationBarrier_25_io_x_c),
    .io_y_ppn(OptimizationBarrier_25_io_y_ppn),
    .io_y_u(OptimizationBarrier_25_io_y_u),
    .io_y_ae(OptimizationBarrier_25_io_y_ae),
    .io_y_sw(OptimizationBarrier_25_io_y_sw),
    .io_y_sx(OptimizationBarrier_25_io_y_sx),
    .io_y_sr(OptimizationBarrier_25_io_y_sr),
    .io_y_pw(OptimizationBarrier_25_io_y_pw),
    .io_y_px(OptimizationBarrier_25_io_y_px),
    .io_y_pr(OptimizationBarrier_25_io_y_pr),
    .io_y_ppp(OptimizationBarrier_25_io_y_ppp),
    .io_y_pal(OptimizationBarrier_25_io_y_pal),
    .io_y_paa(OptimizationBarrier_25_io_y_paa),
    .io_y_eff(OptimizationBarrier_25_io_y_eff),
    .io_y_c(OptimizationBarrier_25_io_y_c),
    .io_covSum(OptimizationBarrier_25_io_covSum),
    .metaAssert(OptimizationBarrier_25_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_26 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_26_io_x_ppn),
    .io_x_u(OptimizationBarrier_26_io_x_u),
    .io_x_ae(OptimizationBarrier_26_io_x_ae),
    .io_x_sw(OptimizationBarrier_26_io_x_sw),
    .io_x_sx(OptimizationBarrier_26_io_x_sx),
    .io_x_sr(OptimizationBarrier_26_io_x_sr),
    .io_x_pw(OptimizationBarrier_26_io_x_pw),
    .io_x_px(OptimizationBarrier_26_io_x_px),
    .io_x_pr(OptimizationBarrier_26_io_x_pr),
    .io_x_ppp(OptimizationBarrier_26_io_x_ppp),
    .io_x_pal(OptimizationBarrier_26_io_x_pal),
    .io_x_paa(OptimizationBarrier_26_io_x_paa),
    .io_x_eff(OptimizationBarrier_26_io_x_eff),
    .io_x_c(OptimizationBarrier_26_io_x_c),
    .io_y_ppn(OptimizationBarrier_26_io_y_ppn),
    .io_y_u(OptimizationBarrier_26_io_y_u),
    .io_y_ae(OptimizationBarrier_26_io_y_ae),
    .io_y_sw(OptimizationBarrier_26_io_y_sw),
    .io_y_sx(OptimizationBarrier_26_io_y_sx),
    .io_y_sr(OptimizationBarrier_26_io_y_sr),
    .io_y_pw(OptimizationBarrier_26_io_y_pw),
    .io_y_px(OptimizationBarrier_26_io_y_px),
    .io_y_pr(OptimizationBarrier_26_io_y_pr),
    .io_y_ppp(OptimizationBarrier_26_io_y_ppp),
    .io_y_pal(OptimizationBarrier_26_io_y_pal),
    .io_y_paa(OptimizationBarrier_26_io_y_paa),
    .io_y_eff(OptimizationBarrier_26_io_y_eff),
    .io_y_c(OptimizationBarrier_26_io_y_c),
    .io_covSum(OptimizationBarrier_26_io_covSum),
    .metaAssert(OptimizationBarrier_26_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_27 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_27_io_x_ppn),
    .io_x_u(OptimizationBarrier_27_io_x_u),
    .io_x_ae(OptimizationBarrier_27_io_x_ae),
    .io_x_sw(OptimizationBarrier_27_io_x_sw),
    .io_x_sx(OptimizationBarrier_27_io_x_sx),
    .io_x_sr(OptimizationBarrier_27_io_x_sr),
    .io_x_pw(OptimizationBarrier_27_io_x_pw),
    .io_x_px(OptimizationBarrier_27_io_x_px),
    .io_x_pr(OptimizationBarrier_27_io_x_pr),
    .io_x_ppp(OptimizationBarrier_27_io_x_ppp),
    .io_x_pal(OptimizationBarrier_27_io_x_pal),
    .io_x_paa(OptimizationBarrier_27_io_x_paa),
    .io_x_eff(OptimizationBarrier_27_io_x_eff),
    .io_x_c(OptimizationBarrier_27_io_x_c),
    .io_y_ppn(OptimizationBarrier_27_io_y_ppn),
    .io_y_u(OptimizationBarrier_27_io_y_u),
    .io_y_ae(OptimizationBarrier_27_io_y_ae),
    .io_y_sw(OptimizationBarrier_27_io_y_sw),
    .io_y_sx(OptimizationBarrier_27_io_y_sx),
    .io_y_sr(OptimizationBarrier_27_io_y_sr),
    .io_y_pw(OptimizationBarrier_27_io_y_pw),
    .io_y_px(OptimizationBarrier_27_io_y_px),
    .io_y_pr(OptimizationBarrier_27_io_y_pr),
    .io_y_ppp(OptimizationBarrier_27_io_y_ppp),
    .io_y_pal(OptimizationBarrier_27_io_y_pal),
    .io_y_paa(OptimizationBarrier_27_io_y_paa),
    .io_y_eff(OptimizationBarrier_27_io_y_eff),
    .io_y_c(OptimizationBarrier_27_io_y_c),
    .io_covSum(OptimizationBarrier_27_io_covSum),
    .metaAssert(OptimizationBarrier_27_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_28 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_28_io_x_ppn),
    .io_x_u(OptimizationBarrier_28_io_x_u),
    .io_x_ae(OptimizationBarrier_28_io_x_ae),
    .io_x_sw(OptimizationBarrier_28_io_x_sw),
    .io_x_sx(OptimizationBarrier_28_io_x_sx),
    .io_x_sr(OptimizationBarrier_28_io_x_sr),
    .io_x_pw(OptimizationBarrier_28_io_x_pw),
    .io_x_px(OptimizationBarrier_28_io_x_px),
    .io_x_pr(OptimizationBarrier_28_io_x_pr),
    .io_x_ppp(OptimizationBarrier_28_io_x_ppp),
    .io_x_pal(OptimizationBarrier_28_io_x_pal),
    .io_x_paa(OptimizationBarrier_28_io_x_paa),
    .io_x_eff(OptimizationBarrier_28_io_x_eff),
    .io_x_c(OptimizationBarrier_28_io_x_c),
    .io_y_ppn(OptimizationBarrier_28_io_y_ppn),
    .io_y_u(OptimizationBarrier_28_io_y_u),
    .io_y_ae(OptimizationBarrier_28_io_y_ae),
    .io_y_sw(OptimizationBarrier_28_io_y_sw),
    .io_y_sx(OptimizationBarrier_28_io_y_sx),
    .io_y_sr(OptimizationBarrier_28_io_y_sr),
    .io_y_pw(OptimizationBarrier_28_io_y_pw),
    .io_y_px(OptimizationBarrier_28_io_y_px),
    .io_y_pr(OptimizationBarrier_28_io_y_pr),
    .io_y_ppp(OptimizationBarrier_28_io_y_ppp),
    .io_y_pal(OptimizationBarrier_28_io_y_pal),
    .io_y_paa(OptimizationBarrier_28_io_y_paa),
    .io_y_eff(OptimizationBarrier_28_io_y_eff),
    .io_y_c(OptimizationBarrier_28_io_y_c),
    .io_covSum(OptimizationBarrier_28_io_covSum),
    .metaAssert(OptimizationBarrier_28_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_29 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_29_io_x_ppn),
    .io_x_u(OptimizationBarrier_29_io_x_u),
    .io_x_ae(OptimizationBarrier_29_io_x_ae),
    .io_x_sw(OptimizationBarrier_29_io_x_sw),
    .io_x_sx(OptimizationBarrier_29_io_x_sx),
    .io_x_sr(OptimizationBarrier_29_io_x_sr),
    .io_x_pw(OptimizationBarrier_29_io_x_pw),
    .io_x_px(OptimizationBarrier_29_io_x_px),
    .io_x_pr(OptimizationBarrier_29_io_x_pr),
    .io_x_ppp(OptimizationBarrier_29_io_x_ppp),
    .io_x_pal(OptimizationBarrier_29_io_x_pal),
    .io_x_paa(OptimizationBarrier_29_io_x_paa),
    .io_x_eff(OptimizationBarrier_29_io_x_eff),
    .io_x_c(OptimizationBarrier_29_io_x_c),
    .io_y_ppn(OptimizationBarrier_29_io_y_ppn),
    .io_y_u(OptimizationBarrier_29_io_y_u),
    .io_y_ae(OptimizationBarrier_29_io_y_ae),
    .io_y_sw(OptimizationBarrier_29_io_y_sw),
    .io_y_sx(OptimizationBarrier_29_io_y_sx),
    .io_y_sr(OptimizationBarrier_29_io_y_sr),
    .io_y_pw(OptimizationBarrier_29_io_y_pw),
    .io_y_px(OptimizationBarrier_29_io_y_px),
    .io_y_pr(OptimizationBarrier_29_io_y_pr),
    .io_y_ppp(OptimizationBarrier_29_io_y_ppp),
    .io_y_pal(OptimizationBarrier_29_io_y_pal),
    .io_y_paa(OptimizationBarrier_29_io_y_paa),
    .io_y_eff(OptimizationBarrier_29_io_y_eff),
    .io_y_c(OptimizationBarrier_29_io_y_c),
    .io_covSum(OptimizationBarrier_29_io_covSum),
    .metaAssert(OptimizationBarrier_29_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_30 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_30_io_x_ppn),
    .io_x_u(OptimizationBarrier_30_io_x_u),
    .io_x_ae(OptimizationBarrier_30_io_x_ae),
    .io_x_sw(OptimizationBarrier_30_io_x_sw),
    .io_x_sx(OptimizationBarrier_30_io_x_sx),
    .io_x_sr(OptimizationBarrier_30_io_x_sr),
    .io_x_pw(OptimizationBarrier_30_io_x_pw),
    .io_x_px(OptimizationBarrier_30_io_x_px),
    .io_x_pr(OptimizationBarrier_30_io_x_pr),
    .io_x_ppp(OptimizationBarrier_30_io_x_ppp),
    .io_x_pal(OptimizationBarrier_30_io_x_pal),
    .io_x_paa(OptimizationBarrier_30_io_x_paa),
    .io_x_eff(OptimizationBarrier_30_io_x_eff),
    .io_x_c(OptimizationBarrier_30_io_x_c),
    .io_y_ppn(OptimizationBarrier_30_io_y_ppn),
    .io_y_u(OptimizationBarrier_30_io_y_u),
    .io_y_ae(OptimizationBarrier_30_io_y_ae),
    .io_y_sw(OptimizationBarrier_30_io_y_sw),
    .io_y_sx(OptimizationBarrier_30_io_y_sx),
    .io_y_sr(OptimizationBarrier_30_io_y_sr),
    .io_y_pw(OptimizationBarrier_30_io_y_pw),
    .io_y_px(OptimizationBarrier_30_io_y_px),
    .io_y_pr(OptimizationBarrier_30_io_y_pr),
    .io_y_ppp(OptimizationBarrier_30_io_y_ppp),
    .io_y_pal(OptimizationBarrier_30_io_y_pal),
    .io_y_paa(OptimizationBarrier_30_io_y_paa),
    .io_y_eff(OptimizationBarrier_30_io_y_eff),
    .io_y_c(OptimizationBarrier_30_io_y_c),
    .io_covSum(OptimizationBarrier_30_io_covSum),
    .metaAssert(OptimizationBarrier_30_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_31 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_31_io_x_ppn),
    .io_x_u(OptimizationBarrier_31_io_x_u),
    .io_x_ae(OptimizationBarrier_31_io_x_ae),
    .io_x_sw(OptimizationBarrier_31_io_x_sw),
    .io_x_sx(OptimizationBarrier_31_io_x_sx),
    .io_x_sr(OptimizationBarrier_31_io_x_sr),
    .io_x_pw(OptimizationBarrier_31_io_x_pw),
    .io_x_px(OptimizationBarrier_31_io_x_px),
    .io_x_pr(OptimizationBarrier_31_io_x_pr),
    .io_x_ppp(OptimizationBarrier_31_io_x_ppp),
    .io_x_pal(OptimizationBarrier_31_io_x_pal),
    .io_x_paa(OptimizationBarrier_31_io_x_paa),
    .io_x_eff(OptimizationBarrier_31_io_x_eff),
    .io_x_c(OptimizationBarrier_31_io_x_c),
    .io_y_ppn(OptimizationBarrier_31_io_y_ppn),
    .io_y_u(OptimizationBarrier_31_io_y_u),
    .io_y_ae(OptimizationBarrier_31_io_y_ae),
    .io_y_sw(OptimizationBarrier_31_io_y_sw),
    .io_y_sx(OptimizationBarrier_31_io_y_sx),
    .io_y_sr(OptimizationBarrier_31_io_y_sr),
    .io_y_pw(OptimizationBarrier_31_io_y_pw),
    .io_y_px(OptimizationBarrier_31_io_y_px),
    .io_y_pr(OptimizationBarrier_31_io_y_pr),
    .io_y_ppp(OptimizationBarrier_31_io_y_ppp),
    .io_y_pal(OptimizationBarrier_31_io_y_pal),
    .io_y_paa(OptimizationBarrier_31_io_y_paa),
    .io_y_eff(OptimizationBarrier_31_io_y_eff),
    .io_y_c(OptimizationBarrier_31_io_y_c),
    .io_covSum(OptimizationBarrier_31_io_covSum),
    .metaAssert(OptimizationBarrier_31_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_32 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_32_io_x_ppn),
    .io_x_u(OptimizationBarrier_32_io_x_u),
    .io_x_ae(OptimizationBarrier_32_io_x_ae),
    .io_x_sw(OptimizationBarrier_32_io_x_sw),
    .io_x_sx(OptimizationBarrier_32_io_x_sx),
    .io_x_sr(OptimizationBarrier_32_io_x_sr),
    .io_x_pw(OptimizationBarrier_32_io_x_pw),
    .io_x_px(OptimizationBarrier_32_io_x_px),
    .io_x_pr(OptimizationBarrier_32_io_x_pr),
    .io_x_ppp(OptimizationBarrier_32_io_x_ppp),
    .io_x_pal(OptimizationBarrier_32_io_x_pal),
    .io_x_paa(OptimizationBarrier_32_io_x_paa),
    .io_x_eff(OptimizationBarrier_32_io_x_eff),
    .io_x_c(OptimizationBarrier_32_io_x_c),
    .io_y_ppn(OptimizationBarrier_32_io_y_ppn),
    .io_y_u(OptimizationBarrier_32_io_y_u),
    .io_y_ae(OptimizationBarrier_32_io_y_ae),
    .io_y_sw(OptimizationBarrier_32_io_y_sw),
    .io_y_sx(OptimizationBarrier_32_io_y_sx),
    .io_y_sr(OptimizationBarrier_32_io_y_sr),
    .io_y_pw(OptimizationBarrier_32_io_y_pw),
    .io_y_px(OptimizationBarrier_32_io_y_px),
    .io_y_pr(OptimizationBarrier_32_io_y_pr),
    .io_y_ppp(OptimizationBarrier_32_io_y_ppp),
    .io_y_pal(OptimizationBarrier_32_io_y_pal),
    .io_y_paa(OptimizationBarrier_32_io_y_paa),
    .io_y_eff(OptimizationBarrier_32_io_y_eff),
    .io_y_c(OptimizationBarrier_32_io_y_c),
    .io_covSum(OptimizationBarrier_32_io_covSum),
    .metaAssert(OptimizationBarrier_32_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_33 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_33_io_x_ppn),
    .io_x_u(OptimizationBarrier_33_io_x_u),
    .io_x_ae(OptimizationBarrier_33_io_x_ae),
    .io_x_sw(OptimizationBarrier_33_io_x_sw),
    .io_x_sx(OptimizationBarrier_33_io_x_sx),
    .io_x_sr(OptimizationBarrier_33_io_x_sr),
    .io_x_pw(OptimizationBarrier_33_io_x_pw),
    .io_x_px(OptimizationBarrier_33_io_x_px),
    .io_x_pr(OptimizationBarrier_33_io_x_pr),
    .io_x_ppp(OptimizationBarrier_33_io_x_ppp),
    .io_x_pal(OptimizationBarrier_33_io_x_pal),
    .io_x_paa(OptimizationBarrier_33_io_x_paa),
    .io_x_eff(OptimizationBarrier_33_io_x_eff),
    .io_x_c(OptimizationBarrier_33_io_x_c),
    .io_y_ppn(OptimizationBarrier_33_io_y_ppn),
    .io_y_u(OptimizationBarrier_33_io_y_u),
    .io_y_ae(OptimizationBarrier_33_io_y_ae),
    .io_y_sw(OptimizationBarrier_33_io_y_sw),
    .io_y_sx(OptimizationBarrier_33_io_y_sx),
    .io_y_sr(OptimizationBarrier_33_io_y_sr),
    .io_y_pw(OptimizationBarrier_33_io_y_pw),
    .io_y_px(OptimizationBarrier_33_io_y_px),
    .io_y_pr(OptimizationBarrier_33_io_y_pr),
    .io_y_ppp(OptimizationBarrier_33_io_y_ppp),
    .io_y_pal(OptimizationBarrier_33_io_y_pal),
    .io_y_paa(OptimizationBarrier_33_io_y_paa),
    .io_y_eff(OptimizationBarrier_33_io_y_eff),
    .io_y_c(OptimizationBarrier_33_io_y_c),
    .io_covSum(OptimizationBarrier_33_io_covSum),
    .metaAssert(OptimizationBarrier_33_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_34 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_34_io_x_ppn),
    .io_x_u(OptimizationBarrier_34_io_x_u),
    .io_x_ae(OptimizationBarrier_34_io_x_ae),
    .io_x_sw(OptimizationBarrier_34_io_x_sw),
    .io_x_sx(OptimizationBarrier_34_io_x_sx),
    .io_x_sr(OptimizationBarrier_34_io_x_sr),
    .io_x_pw(OptimizationBarrier_34_io_x_pw),
    .io_x_px(OptimizationBarrier_34_io_x_px),
    .io_x_pr(OptimizationBarrier_34_io_x_pr),
    .io_x_ppp(OptimizationBarrier_34_io_x_ppp),
    .io_x_pal(OptimizationBarrier_34_io_x_pal),
    .io_x_paa(OptimizationBarrier_34_io_x_paa),
    .io_x_eff(OptimizationBarrier_34_io_x_eff),
    .io_x_c(OptimizationBarrier_34_io_x_c),
    .io_y_ppn(OptimizationBarrier_34_io_y_ppn),
    .io_y_u(OptimizationBarrier_34_io_y_u),
    .io_y_ae(OptimizationBarrier_34_io_y_ae),
    .io_y_sw(OptimizationBarrier_34_io_y_sw),
    .io_y_sx(OptimizationBarrier_34_io_y_sx),
    .io_y_sr(OptimizationBarrier_34_io_y_sr),
    .io_y_pw(OptimizationBarrier_34_io_y_pw),
    .io_y_px(OptimizationBarrier_34_io_y_px),
    .io_y_pr(OptimizationBarrier_34_io_y_pr),
    .io_y_ppp(OptimizationBarrier_34_io_y_ppp),
    .io_y_pal(OptimizationBarrier_34_io_y_pal),
    .io_y_paa(OptimizationBarrier_34_io_y_paa),
    .io_y_eff(OptimizationBarrier_34_io_y_eff),
    .io_y_c(OptimizationBarrier_34_io_y_c),
    .io_covSum(OptimizationBarrier_34_io_covSum),
    .metaAssert(OptimizationBarrier_34_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_35 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_35_io_x_ppn),
    .io_x_u(OptimizationBarrier_35_io_x_u),
    .io_x_ae(OptimizationBarrier_35_io_x_ae),
    .io_x_sw(OptimizationBarrier_35_io_x_sw),
    .io_x_sx(OptimizationBarrier_35_io_x_sx),
    .io_x_sr(OptimizationBarrier_35_io_x_sr),
    .io_x_pw(OptimizationBarrier_35_io_x_pw),
    .io_x_px(OptimizationBarrier_35_io_x_px),
    .io_x_pr(OptimizationBarrier_35_io_x_pr),
    .io_x_ppp(OptimizationBarrier_35_io_x_ppp),
    .io_x_pal(OptimizationBarrier_35_io_x_pal),
    .io_x_paa(OptimizationBarrier_35_io_x_paa),
    .io_x_eff(OptimizationBarrier_35_io_x_eff),
    .io_x_c(OptimizationBarrier_35_io_x_c),
    .io_y_ppn(OptimizationBarrier_35_io_y_ppn),
    .io_y_u(OptimizationBarrier_35_io_y_u),
    .io_y_ae(OptimizationBarrier_35_io_y_ae),
    .io_y_sw(OptimizationBarrier_35_io_y_sw),
    .io_y_sx(OptimizationBarrier_35_io_y_sx),
    .io_y_sr(OptimizationBarrier_35_io_y_sr),
    .io_y_pw(OptimizationBarrier_35_io_y_pw),
    .io_y_px(OptimizationBarrier_35_io_y_px),
    .io_y_pr(OptimizationBarrier_35_io_y_pr),
    .io_y_ppp(OptimizationBarrier_35_io_y_ppp),
    .io_y_pal(OptimizationBarrier_35_io_y_pal),
    .io_y_paa(OptimizationBarrier_35_io_y_paa),
    .io_y_eff(OptimizationBarrier_35_io_y_eff),
    .io_y_c(OptimizationBarrier_35_io_y_c),
    .io_covSum(OptimizationBarrier_35_io_covSum),
    .metaAssert(OptimizationBarrier_35_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_36 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_36_io_x_ppn),
    .io_x_u(OptimizationBarrier_36_io_x_u),
    .io_x_ae(OptimizationBarrier_36_io_x_ae),
    .io_x_sw(OptimizationBarrier_36_io_x_sw),
    .io_x_sx(OptimizationBarrier_36_io_x_sx),
    .io_x_sr(OptimizationBarrier_36_io_x_sr),
    .io_x_pw(OptimizationBarrier_36_io_x_pw),
    .io_x_px(OptimizationBarrier_36_io_x_px),
    .io_x_pr(OptimizationBarrier_36_io_x_pr),
    .io_x_ppp(OptimizationBarrier_36_io_x_ppp),
    .io_x_pal(OptimizationBarrier_36_io_x_pal),
    .io_x_paa(OptimizationBarrier_36_io_x_paa),
    .io_x_eff(OptimizationBarrier_36_io_x_eff),
    .io_x_c(OptimizationBarrier_36_io_x_c),
    .io_y_ppn(OptimizationBarrier_36_io_y_ppn),
    .io_y_u(OptimizationBarrier_36_io_y_u),
    .io_y_ae(OptimizationBarrier_36_io_y_ae),
    .io_y_sw(OptimizationBarrier_36_io_y_sw),
    .io_y_sx(OptimizationBarrier_36_io_y_sx),
    .io_y_sr(OptimizationBarrier_36_io_y_sr),
    .io_y_pw(OptimizationBarrier_36_io_y_pw),
    .io_y_px(OptimizationBarrier_36_io_y_px),
    .io_y_pr(OptimizationBarrier_36_io_y_pr),
    .io_y_ppp(OptimizationBarrier_36_io_y_ppp),
    .io_y_pal(OptimizationBarrier_36_io_y_pal),
    .io_y_paa(OptimizationBarrier_36_io_y_paa),
    .io_y_eff(OptimizationBarrier_36_io_y_eff),
    .io_y_c(OptimizationBarrier_36_io_y_c),
    .io_covSum(OptimizationBarrier_36_io_covSum),
    .metaAssert(OptimizationBarrier_36_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_37 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_37_io_x_ppn),
    .io_x_u(OptimizationBarrier_37_io_x_u),
    .io_x_ae(OptimizationBarrier_37_io_x_ae),
    .io_x_sw(OptimizationBarrier_37_io_x_sw),
    .io_x_sx(OptimizationBarrier_37_io_x_sx),
    .io_x_sr(OptimizationBarrier_37_io_x_sr),
    .io_x_pw(OptimizationBarrier_37_io_x_pw),
    .io_x_px(OptimizationBarrier_37_io_x_px),
    .io_x_pr(OptimizationBarrier_37_io_x_pr),
    .io_x_ppp(OptimizationBarrier_37_io_x_ppp),
    .io_x_pal(OptimizationBarrier_37_io_x_pal),
    .io_x_paa(OptimizationBarrier_37_io_x_paa),
    .io_x_eff(OptimizationBarrier_37_io_x_eff),
    .io_x_c(OptimizationBarrier_37_io_x_c),
    .io_y_ppn(OptimizationBarrier_37_io_y_ppn),
    .io_y_u(OptimizationBarrier_37_io_y_u),
    .io_y_ae(OptimizationBarrier_37_io_y_ae),
    .io_y_sw(OptimizationBarrier_37_io_y_sw),
    .io_y_sx(OptimizationBarrier_37_io_y_sx),
    .io_y_sr(OptimizationBarrier_37_io_y_sr),
    .io_y_pw(OptimizationBarrier_37_io_y_pw),
    .io_y_px(OptimizationBarrier_37_io_y_px),
    .io_y_pr(OptimizationBarrier_37_io_y_pr),
    .io_y_ppp(OptimizationBarrier_37_io_y_ppp),
    .io_y_pal(OptimizationBarrier_37_io_y_pal),
    .io_y_paa(OptimizationBarrier_37_io_y_paa),
    .io_y_eff(OptimizationBarrier_37_io_y_eff),
    .io_y_c(OptimizationBarrier_37_io_y_c),
    .io_covSum(OptimizationBarrier_37_io_covSum),
    .metaAssert(OptimizationBarrier_37_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_38 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_38_io_x_ppn),
    .io_x_u(OptimizationBarrier_38_io_x_u),
    .io_x_ae(OptimizationBarrier_38_io_x_ae),
    .io_x_sw(OptimizationBarrier_38_io_x_sw),
    .io_x_sx(OptimizationBarrier_38_io_x_sx),
    .io_x_sr(OptimizationBarrier_38_io_x_sr),
    .io_x_pw(OptimizationBarrier_38_io_x_pw),
    .io_x_px(OptimizationBarrier_38_io_x_px),
    .io_x_pr(OptimizationBarrier_38_io_x_pr),
    .io_x_ppp(OptimizationBarrier_38_io_x_ppp),
    .io_x_pal(OptimizationBarrier_38_io_x_pal),
    .io_x_paa(OptimizationBarrier_38_io_x_paa),
    .io_x_eff(OptimizationBarrier_38_io_x_eff),
    .io_x_c(OptimizationBarrier_38_io_x_c),
    .io_y_ppn(OptimizationBarrier_38_io_y_ppn),
    .io_y_u(OptimizationBarrier_38_io_y_u),
    .io_y_ae(OptimizationBarrier_38_io_y_ae),
    .io_y_sw(OptimizationBarrier_38_io_y_sw),
    .io_y_sx(OptimizationBarrier_38_io_y_sx),
    .io_y_sr(OptimizationBarrier_38_io_y_sr),
    .io_y_pw(OptimizationBarrier_38_io_y_pw),
    .io_y_px(OptimizationBarrier_38_io_y_px),
    .io_y_pr(OptimizationBarrier_38_io_y_pr),
    .io_y_ppp(OptimizationBarrier_38_io_y_ppp),
    .io_y_pal(OptimizationBarrier_38_io_y_pal),
    .io_y_paa(OptimizationBarrier_38_io_y_paa),
    .io_y_eff(OptimizationBarrier_38_io_y_eff),
    .io_y_c(OptimizationBarrier_38_io_y_c),
    .io_covSum(OptimizationBarrier_38_io_covSum),
    .metaAssert(OptimizationBarrier_38_metaAssert)
  );
  assign priv_s = io_ptw_status_dprv[0]; // @[TLB.scala 177:20]
  assign priv_uses_vm = io_ptw_status_dprv <= 2'h1; // @[TLB.scala 178:27]
  assign _T_2 = io_ptw_ptbr_mode[3] & priv_uses_vm; // @[TLB.scala 179:83]
  assign vm_enabled = _T_2 & ~io_req_bits_passthrough; // @[TLB.scala 179:99]
  assign vpn = io_req_bits_vaddr[38:12]; // @[TLB.scala 182:30]
  assign refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 183:44]
  assign _T_4 = state == 2'h1; // @[package.scala 15:47]
  assign _T_5 = state == 2'h3; // @[package.scala 15:47]
  assign _T_6 = _T_4 | _T_5; // @[package.scala 64:59]
  assign invalidate_refill = _T_6 | io_sfence_valid; // @[TLB.scala 185:88]
  assign _T_27 = special_entry_level < 2'h1; // @[TLB.scala 108:28]
  assign _T_29 = _T_27 ? vpn : 27'h0; // @[TLB.scala 109:28]
  assign _GEN_983 = {{7'd0}, OptimizationBarrier_io_y_ppn}; // @[TLB.scala 109:47]
  assign _T_30 = _T_29 | _GEN_983; // @[TLB.scala 109:47]
  assign _T_33 = special_entry_level < 2'h2; // @[TLB.scala 108:28]
  assign _T_35 = _T_33 ? vpn : 27'h0; // @[TLB.scala 109:28]
  assign _T_36 = _T_35 | _GEN_983; // @[TLB.scala 109:47]
  assign _T_38 = {OptimizationBarrier_io_y_ppn[19:18],_T_30[17:9],_T_36[8:0]}; // @[Cat.scala 29:58]
  assign _T_40 = vm_enabled ? {{8'd0}, _T_38} : io_req_bits_vaddr[39:12]; // @[TLB.scala 187:20]
  assign mpu_ppn = io_ptw_resp_valid ? {{8'd0}, refill_ppn} : _T_40; // @[TLB.scala 186:20]
  assign mpu_physaddr = {mpu_ppn,io_req_bits_vaddr[11:0]}; // @[Cat.scala 29:58]
  assign _T_42 = io_ptw_resp_valid | io_req_bits_passthrough; // @[TLB.scala 189:56]
  assign _T_44 = {io_ptw_status_debug,io_ptw_status_dprv}; // @[Cat.scala 29:58]
  assign mpu_priv = _T_42 ? 3'h1 : _T_44; // @[TLB.scala 189:27]
  assign _T_45 = mpu_physaddr ^ 40'h3000; // @[Parameters.scala 137:31]
  assign _T_46 = {1'b0,$signed(_T_45)}; // @[Parameters.scala 137:49]
  assign _T_48 = $signed(_T_46) & -41'sh1000; // @[Parameters.scala 137:52]
  assign _T_49 = $signed(_T_48) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_50 = mpu_physaddr ^ 40'hc000000; // @[Parameters.scala 137:31]
  assign _T_51 = {1'b0,$signed(_T_50)}; // @[Parameters.scala 137:49]
  assign _T_53 = $signed(_T_51) & -41'sh4000000; // @[Parameters.scala 137:52]
  assign _T_54 = $signed(_T_53) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_55 = mpu_physaddr ^ 40'h2000000; // @[Parameters.scala 137:31]
  assign _T_56 = {1'b0,$signed(_T_55)}; // @[Parameters.scala 137:49]
  assign _T_58 = $signed(_T_56) & -41'sh10000; // @[Parameters.scala 137:52]
  assign _T_59 = $signed(_T_58) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_61 = {1'b0,$signed(mpu_physaddr)}; // @[Parameters.scala 137:49]
  assign _T_63 = $signed(_T_61) & -41'sh1000; // @[Parameters.scala 137:52]
  assign _T_64 = $signed(_T_63) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_65 = mpu_physaddr ^ 40'h10000; // @[Parameters.scala 137:31]
  assign _T_66 = {1'b0,$signed(_T_65)}; // @[Parameters.scala 137:49]
  assign _T_68 = $signed(_T_66) & -41'sh10000; // @[Parameters.scala 137:52]
  assign _T_69 = $signed(_T_68) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_70 = mpu_physaddr ^ 40'h80000000; // @[Parameters.scala 137:31]
  assign _T_71 = {1'b0,$signed(_T_70)}; // @[Parameters.scala 137:49]
  assign _T_73 = $signed(_T_71) & -41'sh10000000; // @[Parameters.scala 137:52]
  assign _T_74 = $signed(_T_73) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_75 = mpu_physaddr ^ 40'h60000000; // @[Parameters.scala 137:31]
  assign _T_76 = {1'b0,$signed(_T_75)}; // @[Parameters.scala 137:49]
  assign _T_78 = $signed(_T_76) & -41'sh20000000; // @[Parameters.scala 137:52]
  assign _T_79 = $signed(_T_78) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_81 = _T_49 | _T_54; // @[TLB.scala 195:67]
  assign _T_82 = _T_81 | _T_59; // @[TLB.scala 195:67]
  assign _T_83 = _T_82 | _T_64; // @[TLB.scala 195:67]
  assign _T_84 = _T_83 | _T_69; // @[TLB.scala 195:67]
  assign _T_85 = _T_84 | _T_74; // @[TLB.scala 195:67]
  assign legal_address = _T_85 | _T_79; // @[TLB.scala 195:67]
  assign _T_94 = $signed(_T_71) & 41'sh80000000; // @[Parameters.scala 137:52]
  assign _T_95 = $signed(_T_94) == 41'sh0; // @[Parameters.scala 137:67]
  assign cacheable = legal_address & _T_95; // @[TLB.scala 197:19]
  assign _T_155 = mpu_physaddr ^ 40'h8000000; // @[Parameters.scala 137:31]
  assign _T_156 = {1'b0,$signed(_T_155)}; // @[Parameters.scala 137:49]
  assign _T_158 = $signed(_T_156) & 41'shc8000000; // @[Parameters.scala 137:52]
  assign _T_159 = $signed(_T_158) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_172 = $signed(_T_61) & 41'shc8010000; // @[Parameters.scala 137:52]
  assign _T_173 = $signed(_T_172) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_180 = _T_173 | _T_159; // @[TLBPermissions.scala 82:66]
  assign _T_193 = mpu_priv <= 3'h3; // @[TLB.scala 200:39]
  assign deny_access_to_debug = _T_193 & _T_64; // @[TLB.scala 200:48]
  assign _T_206 = legal_address & ~deny_access_to_debug; // @[TLB.scala 201:41]
  assign prot_r = _T_206 & pmp_io_r; // @[TLB.scala 201:66]
  assign _T_217 = mpu_physaddr ^ 40'h40000000; // @[Parameters.scala 137:31]
  assign _T_218 = {1'b0,$signed(_T_217)}; // @[Parameters.scala 137:49]
  assign _T_220 = $signed(_T_218) & 41'shc0000000; // @[Parameters.scala 137:52]
  assign _T_221 = $signed(_T_220) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_225 = $signed(_T_71) & 41'shc0000000; // @[Parameters.scala 137:52]
  assign _T_226 = $signed(_T_225) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_228 = _T_180 | _T_221; // @[Parameters.scala 549:89]
  assign _T_229 = _T_228 | _T_226; // @[Parameters.scala 549:89]
  assign _T_239 = legal_address & _T_229; // @[TLB.scala 197:19]
  assign _T_241 = _T_239 & ~deny_access_to_debug; // @[TLB.scala 202:45]
  assign prot_w = _T_241 & pmp_io_w; // @[TLB.scala 202:70]
  assign prot_al = legal_address & _T_180; // @[TLB.scala 197:19]
  assign _T_341 = $signed(_T_61) & 41'shca000000; // @[Parameters.scala 137:52]
  assign _T_342 = $signed(_T_341) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_353 = _T_342 | _T_221; // @[Parameters.scala 549:89]
  assign _T_354 = _T_353 | _T_226; // @[Parameters.scala 549:89]
  assign _T_370 = legal_address & _T_354; // @[TLB.scala 197:19]
  assign _T_372 = _T_370 & ~deny_access_to_debug; // @[TLB.scala 206:40]
  assign prot_x = _T_372 & pmp_io_x; // @[TLB.scala 206:65]
  assign _T_393 = $signed(_T_61) & 41'shca012000; // @[Parameters.scala 137:52]
  assign _T_394 = $signed(_T_393) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_398 = $signed(_T_56) & 41'shca010000; // @[Parameters.scala 137:52]
  assign _T_399 = $signed(_T_398) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_410 = _T_394 | _T_399; // @[Parameters.scala 549:89]
  assign _T_411 = _T_410 | _T_159; // @[Parameters.scala 549:89]
  assign _T_412 = _T_411 | _T_221; // @[Parameters.scala 549:89]
  assign prot_eff = legal_address & _T_412; // @[TLB.scala 197:19]
  assign _T_417 = sectored_entries_0_valid_0 | sectored_entries_0_valid_1; // @[package.scala 64:59]
  assign _T_418 = _T_417 | sectored_entries_0_valid_2; // @[package.scala 64:59]
  assign _T_419 = _T_418 | sectored_entries_0_valid_3; // @[package.scala 64:59]
  assign _T_420 = sectored_entries_0_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_422 = _T_420[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_0 = _T_419 & _T_422; // @[TLB.scala 87:40]
  assign _T_423 = sectored_entries_1_valid_0 | sectored_entries_1_valid_1; // @[package.scala 64:59]
  assign _T_424 = _T_423 | sectored_entries_1_valid_2; // @[package.scala 64:59]
  assign _T_425 = _T_424 | sectored_entries_1_valid_3; // @[package.scala 64:59]
  assign _T_426 = sectored_entries_1_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_428 = _T_426[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_1 = _T_425 & _T_428; // @[TLB.scala 87:40]
  assign _T_429 = sectored_entries_2_valid_0 | sectored_entries_2_valid_1; // @[package.scala 64:59]
  assign _T_430 = _T_429 | sectored_entries_2_valid_2; // @[package.scala 64:59]
  assign _T_431 = _T_430 | sectored_entries_2_valid_3; // @[package.scala 64:59]
  assign _T_432 = sectored_entries_2_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_434 = _T_432[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_2 = _T_431 & _T_434; // @[TLB.scala 87:40]
  assign _T_435 = sectored_entries_3_valid_0 | sectored_entries_3_valid_1; // @[package.scala 64:59]
  assign _T_436 = _T_435 | sectored_entries_3_valid_2; // @[package.scala 64:59]
  assign _T_437 = _T_436 | sectored_entries_3_valid_3; // @[package.scala 64:59]
  assign _T_438 = sectored_entries_3_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_440 = _T_438[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_3 = _T_437 & _T_440; // @[TLB.scala 87:40]
  assign _T_441 = sectored_entries_4_valid_0 | sectored_entries_4_valid_1; // @[package.scala 64:59]
  assign _T_442 = _T_441 | sectored_entries_4_valid_2; // @[package.scala 64:59]
  assign _T_443 = _T_442 | sectored_entries_4_valid_3; // @[package.scala 64:59]
  assign _T_444 = sectored_entries_4_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_446 = _T_444[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_4 = _T_443 & _T_446; // @[TLB.scala 87:40]
  assign _T_447 = sectored_entries_5_valid_0 | sectored_entries_5_valid_1; // @[package.scala 64:59]
  assign _T_448 = _T_447 | sectored_entries_5_valid_2; // @[package.scala 64:59]
  assign _T_449 = _T_448 | sectored_entries_5_valid_3; // @[package.scala 64:59]
  assign _T_450 = sectored_entries_5_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_452 = _T_450[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_5 = _T_449 & _T_452; // @[TLB.scala 87:40]
  assign _T_453 = sectored_entries_6_valid_0 | sectored_entries_6_valid_1; // @[package.scala 64:59]
  assign _T_454 = _T_453 | sectored_entries_6_valid_2; // @[package.scala 64:59]
  assign _T_455 = _T_454 | sectored_entries_6_valid_3; // @[package.scala 64:59]
  assign _T_456 = sectored_entries_6_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_458 = _T_456[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_6 = _T_455 & _T_458; // @[TLB.scala 87:40]
  assign _T_459 = sectored_entries_7_valid_0 | sectored_entries_7_valid_1; // @[package.scala 64:59]
  assign _T_460 = _T_459 | sectored_entries_7_valid_2; // @[package.scala 64:59]
  assign _T_461 = _T_460 | sectored_entries_7_valid_3; // @[package.scala 64:59]
  assign _T_462 = sectored_entries_7_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_464 = _T_462[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_7 = _T_461 & _T_464; // @[TLB.scala 87:40]
  assign _T_469 = superpage_entries_0_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _T_471 = superpage_entries_0_valid_0 & _T_469; // @[TLB.scala 95:29]
  assign _T_472 = superpage_entries_0_level < 2'h1; // @[TLB.scala 94:28]
  assign _T_476 = superpage_entries_0_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _T_477 = _T_472 | _T_476; // @[TLB.scala 95:40]
  assign superpage_hits_0 = _T_471 & _T_477; // @[TLB.scala 95:29]
  assign _T_489 = superpage_entries_1_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _T_491 = superpage_entries_1_valid_0 & _T_489; // @[TLB.scala 95:29]
  assign _T_492 = superpage_entries_1_level < 2'h1; // @[TLB.scala 94:28]
  assign _T_496 = superpage_entries_1_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _T_497 = _T_492 | _T_496; // @[TLB.scala 95:40]
  assign superpage_hits_1 = _T_491 & _T_497; // @[TLB.scala 95:29]
  assign _T_509 = superpage_entries_2_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _T_511 = superpage_entries_2_valid_0 & _T_509; // @[TLB.scala 95:29]
  assign _T_512 = superpage_entries_2_level < 2'h1; // @[TLB.scala 94:28]
  assign _T_516 = superpage_entries_2_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _T_517 = _T_512 | _T_516; // @[TLB.scala 95:40]
  assign superpage_hits_2 = _T_511 & _T_517; // @[TLB.scala 95:29]
  assign _T_529 = superpage_entries_3_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _T_531 = superpage_entries_3_valid_0 & _T_529; // @[TLB.scala 95:29]
  assign _T_532 = superpage_entries_3_level < 2'h1; // @[TLB.scala 94:28]
  assign _T_536 = superpage_entries_3_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _T_537 = _T_532 | _T_536; // @[TLB.scala 95:40]
  assign superpage_hits_3 = _T_531 & _T_537; // @[TLB.scala 95:29]
  assign _GEN_1 = 2'h1 == vpn[1:0] ? sectored_entries_0_valid_1 : sectored_entries_0_valid_0; // @[TLB.scala 100:18]
  assign _GEN_2 = 2'h2 == vpn[1:0] ? sectored_entries_0_valid_2 : _GEN_1; // @[TLB.scala 100:18]
  assign _GEN_3 = 2'h3 == vpn[1:0] ? sectored_entries_0_valid_3 : _GEN_2; // @[TLB.scala 100:18]
  assign _T_549 = _GEN_3 & _T_422; // @[TLB.scala 100:18]
  assign hitsVec_0 = vm_enabled & _T_549; // @[TLB.scala 211:44]
  assign _GEN_5 = 2'h1 == vpn[1:0] ? sectored_entries_1_valid_1 : sectored_entries_1_valid_0; // @[TLB.scala 100:18]
  assign _GEN_6 = 2'h2 == vpn[1:0] ? sectored_entries_1_valid_2 : _GEN_5; // @[TLB.scala 100:18]
  assign _GEN_7 = 2'h3 == vpn[1:0] ? sectored_entries_1_valid_3 : _GEN_6; // @[TLB.scala 100:18]
  assign _T_554 = _GEN_7 & _T_428; // @[TLB.scala 100:18]
  assign hitsVec_1 = vm_enabled & _T_554; // @[TLB.scala 211:44]
  assign _GEN_9 = 2'h1 == vpn[1:0] ? sectored_entries_2_valid_1 : sectored_entries_2_valid_0; // @[TLB.scala 100:18]
  assign _GEN_10 = 2'h2 == vpn[1:0] ? sectored_entries_2_valid_2 : _GEN_9; // @[TLB.scala 100:18]
  assign _GEN_11 = 2'h3 == vpn[1:0] ? sectored_entries_2_valid_3 : _GEN_10; // @[TLB.scala 100:18]
  assign _T_559 = _GEN_11 & _T_434; // @[TLB.scala 100:18]
  assign hitsVec_2 = vm_enabled & _T_559; // @[TLB.scala 211:44]
  assign _GEN_13 = 2'h1 == vpn[1:0] ? sectored_entries_3_valid_1 : sectored_entries_3_valid_0; // @[TLB.scala 100:18]
  assign _GEN_14 = 2'h2 == vpn[1:0] ? sectored_entries_3_valid_2 : _GEN_13; // @[TLB.scala 100:18]
  assign _GEN_15 = 2'h3 == vpn[1:0] ? sectored_entries_3_valid_3 : _GEN_14; // @[TLB.scala 100:18]
  assign _T_564 = _GEN_15 & _T_440; // @[TLB.scala 100:18]
  assign hitsVec_3 = vm_enabled & _T_564; // @[TLB.scala 211:44]
  assign _GEN_17 = 2'h1 == vpn[1:0] ? sectored_entries_4_valid_1 : sectored_entries_4_valid_0; // @[TLB.scala 100:18]
  assign _GEN_18 = 2'h2 == vpn[1:0] ? sectored_entries_4_valid_2 : _GEN_17; // @[TLB.scala 100:18]
  assign _GEN_19 = 2'h3 == vpn[1:0] ? sectored_entries_4_valid_3 : _GEN_18; // @[TLB.scala 100:18]
  assign _T_569 = _GEN_19 & _T_446; // @[TLB.scala 100:18]
  assign hitsVec_4 = vm_enabled & _T_569; // @[TLB.scala 211:44]
  assign _GEN_21 = 2'h1 == vpn[1:0] ? sectored_entries_5_valid_1 : sectored_entries_5_valid_0; // @[TLB.scala 100:18]
  assign _GEN_22 = 2'h2 == vpn[1:0] ? sectored_entries_5_valid_2 : _GEN_21; // @[TLB.scala 100:18]
  assign _GEN_23 = 2'h3 == vpn[1:0] ? sectored_entries_5_valid_3 : _GEN_22; // @[TLB.scala 100:18]
  assign _T_574 = _GEN_23 & _T_452; // @[TLB.scala 100:18]
  assign hitsVec_5 = vm_enabled & _T_574; // @[TLB.scala 211:44]
  assign _GEN_25 = 2'h1 == vpn[1:0] ? sectored_entries_6_valid_1 : sectored_entries_6_valid_0; // @[TLB.scala 100:18]
  assign _GEN_26 = 2'h2 == vpn[1:0] ? sectored_entries_6_valid_2 : _GEN_25; // @[TLB.scala 100:18]
  assign _GEN_27 = 2'h3 == vpn[1:0] ? sectored_entries_6_valid_3 : _GEN_26; // @[TLB.scala 100:18]
  assign _T_579 = _GEN_27 & _T_458; // @[TLB.scala 100:18]
  assign hitsVec_6 = vm_enabled & _T_579; // @[TLB.scala 211:44]
  assign _GEN_29 = 2'h1 == vpn[1:0] ? sectored_entries_7_valid_1 : sectored_entries_7_valid_0; // @[TLB.scala 100:18]
  assign _GEN_30 = 2'h2 == vpn[1:0] ? sectored_entries_7_valid_2 : _GEN_29; // @[TLB.scala 100:18]
  assign _GEN_31 = 2'h3 == vpn[1:0] ? sectored_entries_7_valid_3 : _GEN_30; // @[TLB.scala 100:18]
  assign _T_584 = _GEN_31 & _T_464; // @[TLB.scala 100:18]
  assign hitsVec_7 = vm_enabled & _T_584; // @[TLB.scala 211:44]
  assign hitsVec_8 = vm_enabled & superpage_hits_0; // @[TLB.scala 211:44]
  assign hitsVec_9 = vm_enabled & superpage_hits_1; // @[TLB.scala 211:44]
  assign hitsVec_10 = vm_enabled & superpage_hits_2; // @[TLB.scala 211:44]
  assign hitsVec_11 = vm_enabled & superpage_hits_3; // @[TLB.scala 211:44]
  assign _T_673 = special_entry_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _T_675 = special_entry_valid_0 & _T_673; // @[TLB.scala 95:29]
  assign _T_680 = special_entry_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _T_681 = _T_27 | _T_680; // @[TLB.scala 95:40]
  assign _T_682 = _T_675 & _T_681; // @[TLB.scala 95:29]
  assign _T_687 = special_entry_tag[8:0] == vpn[8:0]; // @[TLB.scala 95:77]
  assign _T_688 = _T_33 | _T_687; // @[TLB.scala 95:40]
  assign _T_689 = _T_682 & _T_688; // @[TLB.scala 95:29]
  assign hitsVec_12 = vm_enabled & _T_689; // @[TLB.scala 211:44]
  assign _T_694 = {hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[Cat.scala 29:58]
  assign real_hits = {hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_694}; // @[Cat.scala 29:58]
  assign hits = {~vm_enabled,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_694}; // @[Cat.scala 29:58]
  assign _GEN_33 = 2'h1 == vpn[1:0] ? sectored_entries_0_data_1 : sectored_entries_0_data_0;
  assign _GEN_34 = 2'h2 == vpn[1:0] ? sectored_entries_0_data_2 : _GEN_33;
  assign _GEN_35 = 2'h3 == vpn[1:0] ? sectored_entries_0_data_3 : _GEN_34;
  assign _GEN_37 = 2'h1 == vpn[1:0] ? sectored_entries_1_data_1 : sectored_entries_1_data_0;
  assign _GEN_38 = 2'h2 == vpn[1:0] ? sectored_entries_1_data_2 : _GEN_37;
  assign _GEN_39 = 2'h3 == vpn[1:0] ? sectored_entries_1_data_3 : _GEN_38;
  assign _GEN_41 = 2'h1 == vpn[1:0] ? sectored_entries_2_data_1 : sectored_entries_2_data_0;
  assign _GEN_42 = 2'h2 == vpn[1:0] ? sectored_entries_2_data_2 : _GEN_41;
  assign _GEN_43 = 2'h3 == vpn[1:0] ? sectored_entries_2_data_3 : _GEN_42;
  assign _GEN_45 = 2'h1 == vpn[1:0] ? sectored_entries_3_data_1 : sectored_entries_3_data_0;
  assign _GEN_46 = 2'h2 == vpn[1:0] ? sectored_entries_3_data_2 : _GEN_45;
  assign _GEN_47 = 2'h3 == vpn[1:0] ? sectored_entries_3_data_3 : _GEN_46;
  assign _GEN_49 = 2'h1 == vpn[1:0] ? sectored_entries_4_data_1 : sectored_entries_4_data_0;
  assign _GEN_50 = 2'h2 == vpn[1:0] ? sectored_entries_4_data_2 : _GEN_49;
  assign _GEN_51 = 2'h3 == vpn[1:0] ? sectored_entries_4_data_3 : _GEN_50;
  assign _GEN_53 = 2'h1 == vpn[1:0] ? sectored_entries_5_data_1 : sectored_entries_5_data_0;
  assign _GEN_54 = 2'h2 == vpn[1:0] ? sectored_entries_5_data_2 : _GEN_53;
  assign _GEN_55 = 2'h3 == vpn[1:0] ? sectored_entries_5_data_3 : _GEN_54;
  assign _GEN_57 = 2'h1 == vpn[1:0] ? sectored_entries_6_data_1 : sectored_entries_6_data_0;
  assign _GEN_58 = 2'h2 == vpn[1:0] ? sectored_entries_6_data_2 : _GEN_57;
  assign _GEN_59 = 2'h3 == vpn[1:0] ? sectored_entries_6_data_3 : _GEN_58;
  assign _GEN_61 = 2'h1 == vpn[1:0] ? sectored_entries_7_data_1 : sectored_entries_7_data_0;
  assign _GEN_62 = 2'h2 == vpn[1:0] ? sectored_entries_7_data_2 : _GEN_61;
  assign _GEN_63 = 2'h3 == vpn[1:0] ? sectored_entries_7_data_3 : _GEN_62;
  assign _T_876 = _T_472 ? vpn : 27'h0; // @[TLB.scala 109:28]
  assign _GEN_985 = {{7'd0}, OptimizationBarrier_9_io_y_ppn}; // @[TLB.scala 109:47]
  assign _T_877 = _T_876 | _GEN_985; // @[TLB.scala 109:47]
  assign _T_883 = vpn | _GEN_985; // @[TLB.scala 109:47]
  assign _T_885 = {OptimizationBarrier_9_io_y_ppn[19:18],_T_877[17:9],_T_883[8:0]}; // @[Cat.scala 29:58]
  assign _T_907 = _T_492 ? vpn : 27'h0; // @[TLB.scala 109:28]
  assign _GEN_987 = {{7'd0}, OptimizationBarrier_10_io_y_ppn}; // @[TLB.scala 109:47]
  assign _T_908 = _T_907 | _GEN_987; // @[TLB.scala 109:47]
  assign _T_914 = vpn | _GEN_987; // @[TLB.scala 109:47]
  assign _T_916 = {OptimizationBarrier_10_io_y_ppn[19:18],_T_908[17:9],_T_914[8:0]}; // @[Cat.scala 29:58]
  assign _T_938 = _T_512 ? vpn : 27'h0; // @[TLB.scala 109:28]
  assign _GEN_989 = {{7'd0}, OptimizationBarrier_11_io_y_ppn}; // @[TLB.scala 109:47]
  assign _T_939 = _T_938 | _GEN_989; // @[TLB.scala 109:47]
  assign _T_945 = vpn | _GEN_989; // @[TLB.scala 109:47]
  assign _T_947 = {OptimizationBarrier_11_io_y_ppn[19:18],_T_939[17:9],_T_945[8:0]}; // @[Cat.scala 29:58]
  assign _T_969 = _T_532 ? vpn : 27'h0; // @[TLB.scala 109:28]
  assign _GEN_991 = {{7'd0}, OptimizationBarrier_12_io_y_ppn}; // @[TLB.scala 109:47]
  assign _T_970 = _T_969 | _GEN_991; // @[TLB.scala 109:47]
  assign _T_976 = vpn | _GEN_991; // @[TLB.scala 109:47]
  assign _T_978 = {OptimizationBarrier_12_io_y_ppn[19:18],_T_970[17:9],_T_976[8:0]}; // @[Cat.scala 29:58]
  assign _GEN_993 = {{7'd0}, OptimizationBarrier_13_io_y_ppn}; // @[TLB.scala 109:47]
  assign _T_1001 = _T_29 | _GEN_993; // @[TLB.scala 109:47]
  assign _T_1007 = _T_35 | _GEN_993; // @[TLB.scala 109:47]
  assign _T_1009 = {OptimizationBarrier_13_io_y_ppn[19:18],_T_1001[17:9],_T_1007[8:0]}; // @[Cat.scala 29:58]
  assign _T_1011 = hitsVec_0 ? OptimizationBarrier_1_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1012 = hitsVec_1 ? OptimizationBarrier_2_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1013 = hitsVec_2 ? OptimizationBarrier_3_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1014 = hitsVec_3 ? OptimizationBarrier_4_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1015 = hitsVec_4 ? OptimizationBarrier_5_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1016 = hitsVec_5 ? OptimizationBarrier_6_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1017 = hitsVec_6 ? OptimizationBarrier_7_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1018 = hitsVec_7 ? OptimizationBarrier_8_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1019 = hitsVec_8 ? _T_885 : 20'h0; // @[Mux.scala 27:72]
  assign _T_1020 = hitsVec_9 ? _T_916 : 20'h0; // @[Mux.scala 27:72]
  assign _T_1021 = hitsVec_10 ? _T_947 : 20'h0; // @[Mux.scala 27:72]
  assign _T_1022 = hitsVec_11 ? _T_978 : 20'h0; // @[Mux.scala 27:72]
  assign _T_1023 = hitsVec_12 ? _T_1009 : 20'h0; // @[Mux.scala 27:72]
  assign _T_1024 = vm_enabled ? 20'h0 : vpn[19:0]; // @[Mux.scala 27:72]
  assign _T_1025 = _T_1011 | _T_1012; // @[Mux.scala 27:72]
  assign _T_1026 = _T_1025 | _T_1013; // @[Mux.scala 27:72]
  assign _T_1027 = _T_1026 | _T_1014; // @[Mux.scala 27:72]
  assign _T_1028 = _T_1027 | _T_1015; // @[Mux.scala 27:72]
  assign _T_1029 = _T_1028 | _T_1016; // @[Mux.scala 27:72]
  assign _T_1030 = _T_1029 | _T_1017; // @[Mux.scala 27:72]
  assign _T_1031 = _T_1030 | _T_1018; // @[Mux.scala 27:72]
  assign _T_1032 = _T_1031 | _T_1019; // @[Mux.scala 27:72]
  assign _T_1033 = _T_1032 | _T_1020; // @[Mux.scala 27:72]
  assign _T_1034 = _T_1033 | _T_1021; // @[Mux.scala 27:72]
  assign _T_1035 = _T_1034 | _T_1022; // @[Mux.scala 27:72]
  assign _T_1036 = _T_1035 | _T_1023; // @[Mux.scala 27:72]
  assign ppn = _T_1036 | _T_1024; // @[Mux.scala 27:72]
  assign _T_1039 = io_ptw_resp_bits_pte_g & io_ptw_resp_bits_pte_v; // @[TLB.scala 223:25]
  assign _T_1041 = io_ptw_resp_bits_pte_x & ~io_ptw_resp_bits_pte_w; // @[PTW.scala 69:44]
  assign _T_1042 = io_ptw_resp_bits_pte_r | _T_1041; // @[PTW.scala 69:38]
  assign _T_1043 = io_ptw_resp_bits_pte_v & _T_1042; // @[PTW.scala 69:32]
  assign _T_1044 = _T_1043 & io_ptw_resp_bits_pte_a; // @[PTW.scala 69:52]
  assign _T_1045 = _T_1044 & io_ptw_resp_bits_pte_r; // @[PTW.scala 73:35]
  assign _T_1051 = _T_1044 & io_ptw_resp_bits_pte_w; // @[PTW.scala 74:35]
  assign _T_1052 = _T_1051 & io_ptw_resp_bits_pte_d; // @[PTW.scala 74:40]
  assign _T_1058 = _T_1044 & io_ptw_resp_bits_pte_x; // @[PTW.scala 75:35]
  assign _T_1068 = {prot_x,prot_r,_T_239,prot_al,prot_al,prot_eff,cacheable,1'h0}; // @[TLB.scala 123:24]
  assign _T_1076 = {refill_ppn,io_ptw_resp_bits_pte_u,_T_1039,io_ptw_resp_bits_ae,_T_1052,_T_1058,_T_1045,prot_w,_T_1068}; // @[TLB.scala 123:24]
  assign _GEN_64 = invalidate_refill ? 1'h0 : 1'h1; // @[TLB.scala 240:34]
  assign _T_1077 = io_ptw_resp_bits_level < 2'h2; // @[TLB.scala 242:40]
  assign _T_1078 = r_superpage_repl_addr == 2'h0; // @[TLB.scala 243:82]
  assign _GEN_67 = _T_1078 ? _GEN_64 : superpage_entries_0_valid_0; // @[TLB.scala 243:89]
  assign _T_1095 = r_superpage_repl_addr == 2'h1; // @[TLB.scala 243:82]
  assign _GEN_71 = _T_1095 ? _GEN_64 : superpage_entries_1_valid_0; // @[TLB.scala 243:89]
  assign _T_1112 = r_superpage_repl_addr == 2'h2; // @[TLB.scala 243:82]
  assign _GEN_75 = _T_1112 ? _GEN_64 : superpage_entries_2_valid_0; // @[TLB.scala 243:89]
  assign _T_1129 = r_superpage_repl_addr == 2'h3; // @[TLB.scala 243:82]
  assign _GEN_79 = _T_1129 ? _GEN_64 : superpage_entries_3_valid_0; // @[TLB.scala 243:89]
  assign _T_1146 = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; // @[TLB.scala 248:22]
  assign _T_1147 = _T_1146 == 3'h0; // @[TLB.scala 249:65]
  assign _GEN_81 = r_sectored_hit ? sectored_entries_0_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_82 = r_sectored_hit ? sectored_entries_0_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_83 = r_sectored_hit ? sectored_entries_0_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_84 = r_sectored_hit ? sectored_entries_0_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_995 = 2'h0 == r_refill_tag[1:0]; // @[TLB.scala 122:16]
  assign _GEN_85 = _GEN_995 | _GEN_81; // @[TLB.scala 122:16]
  assign _GEN_996 = 2'h1 == r_refill_tag[1:0]; // @[TLB.scala 122:16]
  assign _GEN_86 = _GEN_996 | _GEN_82; // @[TLB.scala 122:16]
  assign _GEN_997 = 2'h2 == r_refill_tag[1:0]; // @[TLB.scala 122:16]
  assign _GEN_87 = _GEN_997 | _GEN_83; // @[TLB.scala 122:16]
  assign _GEN_998 = 2'h3 == r_refill_tag[1:0]; // @[TLB.scala 122:16]
  assign _GEN_88 = _GEN_998 | _GEN_84; // @[TLB.scala 122:16]
  assign _GEN_93 = invalidate_refill ? 1'h0 : _GEN_85; // @[TLB.scala 252:34]
  assign _GEN_94 = invalidate_refill ? 1'h0 : _GEN_86; // @[TLB.scala 252:34]
  assign _GEN_95 = invalidate_refill ? 1'h0 : _GEN_87; // @[TLB.scala 252:34]
  assign _GEN_96 = invalidate_refill ? 1'h0 : _GEN_88; // @[TLB.scala 252:34]
  assign _GEN_97 = _T_1147 ? _GEN_93 : sectored_entries_0_valid_0; // @[TLB.scala 249:72]
  assign _GEN_98 = _T_1147 ? _GEN_94 : sectored_entries_0_valid_1; // @[TLB.scala 249:72]
  assign _GEN_99 = _T_1147 ? _GEN_95 : sectored_entries_0_valid_2; // @[TLB.scala 249:72]
  assign _GEN_100 = _T_1147 ? _GEN_96 : sectored_entries_0_valid_3; // @[TLB.scala 249:72]
  assign _T_1165 = _T_1146 == 3'h1; // @[TLB.scala 249:65]
  assign _GEN_107 = r_sectored_hit ? sectored_entries_1_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_108 = r_sectored_hit ? sectored_entries_1_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_109 = r_sectored_hit ? sectored_entries_1_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_110 = r_sectored_hit ? sectored_entries_1_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_111 = _GEN_995 | _GEN_107; // @[TLB.scala 122:16]
  assign _GEN_112 = _GEN_996 | _GEN_108; // @[TLB.scala 122:16]
  assign _GEN_113 = _GEN_997 | _GEN_109; // @[TLB.scala 122:16]
  assign _GEN_114 = _GEN_998 | _GEN_110; // @[TLB.scala 122:16]
  assign _GEN_119 = invalidate_refill ? 1'h0 : _GEN_111; // @[TLB.scala 252:34]
  assign _GEN_120 = invalidate_refill ? 1'h0 : _GEN_112; // @[TLB.scala 252:34]
  assign _GEN_121 = invalidate_refill ? 1'h0 : _GEN_113; // @[TLB.scala 252:34]
  assign _GEN_122 = invalidate_refill ? 1'h0 : _GEN_114; // @[TLB.scala 252:34]
  assign _GEN_123 = _T_1165 ? _GEN_119 : sectored_entries_1_valid_0; // @[TLB.scala 249:72]
  assign _GEN_124 = _T_1165 ? _GEN_120 : sectored_entries_1_valid_1; // @[TLB.scala 249:72]
  assign _GEN_125 = _T_1165 ? _GEN_121 : sectored_entries_1_valid_2; // @[TLB.scala 249:72]
  assign _GEN_126 = _T_1165 ? _GEN_122 : sectored_entries_1_valid_3; // @[TLB.scala 249:72]
  assign _T_1183 = _T_1146 == 3'h2; // @[TLB.scala 249:65]
  assign _GEN_133 = r_sectored_hit ? sectored_entries_2_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_134 = r_sectored_hit ? sectored_entries_2_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_135 = r_sectored_hit ? sectored_entries_2_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_136 = r_sectored_hit ? sectored_entries_2_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_137 = _GEN_995 | _GEN_133; // @[TLB.scala 122:16]
  assign _GEN_138 = _GEN_996 | _GEN_134; // @[TLB.scala 122:16]
  assign _GEN_139 = _GEN_997 | _GEN_135; // @[TLB.scala 122:16]
  assign _GEN_140 = _GEN_998 | _GEN_136; // @[TLB.scala 122:16]
  assign _GEN_145 = invalidate_refill ? 1'h0 : _GEN_137; // @[TLB.scala 252:34]
  assign _GEN_146 = invalidate_refill ? 1'h0 : _GEN_138; // @[TLB.scala 252:34]
  assign _GEN_147 = invalidate_refill ? 1'h0 : _GEN_139; // @[TLB.scala 252:34]
  assign _GEN_148 = invalidate_refill ? 1'h0 : _GEN_140; // @[TLB.scala 252:34]
  assign _GEN_149 = _T_1183 ? _GEN_145 : sectored_entries_2_valid_0; // @[TLB.scala 249:72]
  assign _GEN_150 = _T_1183 ? _GEN_146 : sectored_entries_2_valid_1; // @[TLB.scala 249:72]
  assign _GEN_151 = _T_1183 ? _GEN_147 : sectored_entries_2_valid_2; // @[TLB.scala 249:72]
  assign _GEN_152 = _T_1183 ? _GEN_148 : sectored_entries_2_valid_3; // @[TLB.scala 249:72]
  assign _T_1201 = _T_1146 == 3'h3; // @[TLB.scala 249:65]
  assign _GEN_159 = r_sectored_hit ? sectored_entries_3_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_160 = r_sectored_hit ? sectored_entries_3_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_161 = r_sectored_hit ? sectored_entries_3_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_162 = r_sectored_hit ? sectored_entries_3_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_163 = _GEN_995 | _GEN_159; // @[TLB.scala 122:16]
  assign _GEN_164 = _GEN_996 | _GEN_160; // @[TLB.scala 122:16]
  assign _GEN_165 = _GEN_997 | _GEN_161; // @[TLB.scala 122:16]
  assign _GEN_166 = _GEN_998 | _GEN_162; // @[TLB.scala 122:16]
  assign _GEN_171 = invalidate_refill ? 1'h0 : _GEN_163; // @[TLB.scala 252:34]
  assign _GEN_172 = invalidate_refill ? 1'h0 : _GEN_164; // @[TLB.scala 252:34]
  assign _GEN_173 = invalidate_refill ? 1'h0 : _GEN_165; // @[TLB.scala 252:34]
  assign _GEN_174 = invalidate_refill ? 1'h0 : _GEN_166; // @[TLB.scala 252:34]
  assign _GEN_175 = _T_1201 ? _GEN_171 : sectored_entries_3_valid_0; // @[TLB.scala 249:72]
  assign _GEN_176 = _T_1201 ? _GEN_172 : sectored_entries_3_valid_1; // @[TLB.scala 249:72]
  assign _GEN_177 = _T_1201 ? _GEN_173 : sectored_entries_3_valid_2; // @[TLB.scala 249:72]
  assign _GEN_178 = _T_1201 ? _GEN_174 : sectored_entries_3_valid_3; // @[TLB.scala 249:72]
  assign _T_1219 = _T_1146 == 3'h4; // @[TLB.scala 249:65]
  assign _GEN_185 = r_sectored_hit ? sectored_entries_4_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_186 = r_sectored_hit ? sectored_entries_4_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_187 = r_sectored_hit ? sectored_entries_4_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_188 = r_sectored_hit ? sectored_entries_4_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_189 = _GEN_995 | _GEN_185; // @[TLB.scala 122:16]
  assign _GEN_190 = _GEN_996 | _GEN_186; // @[TLB.scala 122:16]
  assign _GEN_191 = _GEN_997 | _GEN_187; // @[TLB.scala 122:16]
  assign _GEN_192 = _GEN_998 | _GEN_188; // @[TLB.scala 122:16]
  assign _GEN_197 = invalidate_refill ? 1'h0 : _GEN_189; // @[TLB.scala 252:34]
  assign _GEN_198 = invalidate_refill ? 1'h0 : _GEN_190; // @[TLB.scala 252:34]
  assign _GEN_199 = invalidate_refill ? 1'h0 : _GEN_191; // @[TLB.scala 252:34]
  assign _GEN_200 = invalidate_refill ? 1'h0 : _GEN_192; // @[TLB.scala 252:34]
  assign _GEN_201 = _T_1219 ? _GEN_197 : sectored_entries_4_valid_0; // @[TLB.scala 249:72]
  assign _GEN_202 = _T_1219 ? _GEN_198 : sectored_entries_4_valid_1; // @[TLB.scala 249:72]
  assign _GEN_203 = _T_1219 ? _GEN_199 : sectored_entries_4_valid_2; // @[TLB.scala 249:72]
  assign _GEN_204 = _T_1219 ? _GEN_200 : sectored_entries_4_valid_3; // @[TLB.scala 249:72]
  assign _T_1237 = _T_1146 == 3'h5; // @[TLB.scala 249:65]
  assign _GEN_211 = r_sectored_hit ? sectored_entries_5_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_212 = r_sectored_hit ? sectored_entries_5_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_213 = r_sectored_hit ? sectored_entries_5_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_214 = r_sectored_hit ? sectored_entries_5_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_215 = _GEN_995 | _GEN_211; // @[TLB.scala 122:16]
  assign _GEN_216 = _GEN_996 | _GEN_212; // @[TLB.scala 122:16]
  assign _GEN_217 = _GEN_997 | _GEN_213; // @[TLB.scala 122:16]
  assign _GEN_218 = _GEN_998 | _GEN_214; // @[TLB.scala 122:16]
  assign _GEN_223 = invalidate_refill ? 1'h0 : _GEN_215; // @[TLB.scala 252:34]
  assign _GEN_224 = invalidate_refill ? 1'h0 : _GEN_216; // @[TLB.scala 252:34]
  assign _GEN_225 = invalidate_refill ? 1'h0 : _GEN_217; // @[TLB.scala 252:34]
  assign _GEN_226 = invalidate_refill ? 1'h0 : _GEN_218; // @[TLB.scala 252:34]
  assign _GEN_227 = _T_1237 ? _GEN_223 : sectored_entries_5_valid_0; // @[TLB.scala 249:72]
  assign _GEN_228 = _T_1237 ? _GEN_224 : sectored_entries_5_valid_1; // @[TLB.scala 249:72]
  assign _GEN_229 = _T_1237 ? _GEN_225 : sectored_entries_5_valid_2; // @[TLB.scala 249:72]
  assign _GEN_230 = _T_1237 ? _GEN_226 : sectored_entries_5_valid_3; // @[TLB.scala 249:72]
  assign _T_1255 = _T_1146 == 3'h6; // @[TLB.scala 249:65]
  assign _GEN_237 = r_sectored_hit ? sectored_entries_6_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_238 = r_sectored_hit ? sectored_entries_6_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_239 = r_sectored_hit ? sectored_entries_6_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_240 = r_sectored_hit ? sectored_entries_6_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_241 = _GEN_995 | _GEN_237; // @[TLB.scala 122:16]
  assign _GEN_242 = _GEN_996 | _GEN_238; // @[TLB.scala 122:16]
  assign _GEN_243 = _GEN_997 | _GEN_239; // @[TLB.scala 122:16]
  assign _GEN_244 = _GEN_998 | _GEN_240; // @[TLB.scala 122:16]
  assign _GEN_249 = invalidate_refill ? 1'h0 : _GEN_241; // @[TLB.scala 252:34]
  assign _GEN_250 = invalidate_refill ? 1'h0 : _GEN_242; // @[TLB.scala 252:34]
  assign _GEN_251 = invalidate_refill ? 1'h0 : _GEN_243; // @[TLB.scala 252:34]
  assign _GEN_252 = invalidate_refill ? 1'h0 : _GEN_244; // @[TLB.scala 252:34]
  assign _GEN_253 = _T_1255 ? _GEN_249 : sectored_entries_6_valid_0; // @[TLB.scala 249:72]
  assign _GEN_254 = _T_1255 ? _GEN_250 : sectored_entries_6_valid_1; // @[TLB.scala 249:72]
  assign _GEN_255 = _T_1255 ? _GEN_251 : sectored_entries_6_valid_2; // @[TLB.scala 249:72]
  assign _GEN_256 = _T_1255 ? _GEN_252 : sectored_entries_6_valid_3; // @[TLB.scala 249:72]
  assign _T_1273 = _T_1146 == 3'h7; // @[TLB.scala 249:65]
  assign _GEN_263 = r_sectored_hit ? sectored_entries_7_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_264 = r_sectored_hit ? sectored_entries_7_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_265 = r_sectored_hit ? sectored_entries_7_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_266 = r_sectored_hit ? sectored_entries_7_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_267 = _GEN_995 | _GEN_263; // @[TLB.scala 122:16]
  assign _GEN_268 = _GEN_996 | _GEN_264; // @[TLB.scala 122:16]
  assign _GEN_269 = _GEN_997 | _GEN_265; // @[TLB.scala 122:16]
  assign _GEN_270 = _GEN_998 | _GEN_266; // @[TLB.scala 122:16]
  assign _GEN_275 = invalidate_refill ? 1'h0 : _GEN_267; // @[TLB.scala 252:34]
  assign _GEN_276 = invalidate_refill ? 1'h0 : _GEN_268; // @[TLB.scala 252:34]
  assign _GEN_277 = invalidate_refill ? 1'h0 : _GEN_269; // @[TLB.scala 252:34]
  assign _GEN_278 = invalidate_refill ? 1'h0 : _GEN_270; // @[TLB.scala 252:34]
  assign _GEN_279 = _T_1273 ? _GEN_275 : sectored_entries_7_valid_0; // @[TLB.scala 249:72]
  assign _GEN_280 = _T_1273 ? _GEN_276 : sectored_entries_7_valid_1; // @[TLB.scala 249:72]
  assign _GEN_281 = _T_1273 ? _GEN_277 : sectored_entries_7_valid_2; // @[TLB.scala 249:72]
  assign _GEN_282 = _T_1273 ? _GEN_278 : sectored_entries_7_valid_3; // @[TLB.scala 249:72]
  assign _GEN_291 = _T_1077 ? _GEN_67 : superpage_entries_0_valid_0; // @[TLB.scala 242:54]
  assign _GEN_295 = _T_1077 ? _GEN_71 : superpage_entries_1_valid_0; // @[TLB.scala 242:54]
  assign _GEN_299 = _T_1077 ? _GEN_75 : superpage_entries_2_valid_0; // @[TLB.scala 242:54]
  assign _GEN_303 = _T_1077 ? _GEN_79 : superpage_entries_3_valid_0; // @[TLB.scala 242:54]
  assign _GEN_305 = _T_1077 ? sectored_entries_0_valid_0 : _GEN_97; // @[TLB.scala 242:54]
  assign _GEN_306 = _T_1077 ? sectored_entries_0_valid_1 : _GEN_98; // @[TLB.scala 242:54]
  assign _GEN_307 = _T_1077 ? sectored_entries_0_valid_2 : _GEN_99; // @[TLB.scala 242:54]
  assign _GEN_308 = _T_1077 ? sectored_entries_0_valid_3 : _GEN_100; // @[TLB.scala 242:54]
  assign _GEN_315 = _T_1077 ? sectored_entries_1_valid_0 : _GEN_123; // @[TLB.scala 242:54]
  assign _GEN_316 = _T_1077 ? sectored_entries_1_valid_1 : _GEN_124; // @[TLB.scala 242:54]
  assign _GEN_317 = _T_1077 ? sectored_entries_1_valid_2 : _GEN_125; // @[TLB.scala 242:54]
  assign _GEN_318 = _T_1077 ? sectored_entries_1_valid_3 : _GEN_126; // @[TLB.scala 242:54]
  assign _GEN_325 = _T_1077 ? sectored_entries_2_valid_0 : _GEN_149; // @[TLB.scala 242:54]
  assign _GEN_326 = _T_1077 ? sectored_entries_2_valid_1 : _GEN_150; // @[TLB.scala 242:54]
  assign _GEN_327 = _T_1077 ? sectored_entries_2_valid_2 : _GEN_151; // @[TLB.scala 242:54]
  assign _GEN_328 = _T_1077 ? sectored_entries_2_valid_3 : _GEN_152; // @[TLB.scala 242:54]
  assign _GEN_335 = _T_1077 ? sectored_entries_3_valid_0 : _GEN_175; // @[TLB.scala 242:54]
  assign _GEN_336 = _T_1077 ? sectored_entries_3_valid_1 : _GEN_176; // @[TLB.scala 242:54]
  assign _GEN_337 = _T_1077 ? sectored_entries_3_valid_2 : _GEN_177; // @[TLB.scala 242:54]
  assign _GEN_338 = _T_1077 ? sectored_entries_3_valid_3 : _GEN_178; // @[TLB.scala 242:54]
  assign _GEN_345 = _T_1077 ? sectored_entries_4_valid_0 : _GEN_201; // @[TLB.scala 242:54]
  assign _GEN_346 = _T_1077 ? sectored_entries_4_valid_1 : _GEN_202; // @[TLB.scala 242:54]
  assign _GEN_347 = _T_1077 ? sectored_entries_4_valid_2 : _GEN_203; // @[TLB.scala 242:54]
  assign _GEN_348 = _T_1077 ? sectored_entries_4_valid_3 : _GEN_204; // @[TLB.scala 242:54]
  assign _GEN_355 = _T_1077 ? sectored_entries_5_valid_0 : _GEN_227; // @[TLB.scala 242:54]
  assign _GEN_356 = _T_1077 ? sectored_entries_5_valid_1 : _GEN_228; // @[TLB.scala 242:54]
  assign _GEN_357 = _T_1077 ? sectored_entries_5_valid_2 : _GEN_229; // @[TLB.scala 242:54]
  assign _GEN_358 = _T_1077 ? sectored_entries_5_valid_3 : _GEN_230; // @[TLB.scala 242:54]
  assign _GEN_365 = _T_1077 ? sectored_entries_6_valid_0 : _GEN_253; // @[TLB.scala 242:54]
  assign _GEN_366 = _T_1077 ? sectored_entries_6_valid_1 : _GEN_254; // @[TLB.scala 242:54]
  assign _GEN_367 = _T_1077 ? sectored_entries_6_valid_2 : _GEN_255; // @[TLB.scala 242:54]
  assign _GEN_368 = _T_1077 ? sectored_entries_6_valid_3 : _GEN_256; // @[TLB.scala 242:54]
  assign _GEN_375 = _T_1077 ? sectored_entries_7_valid_0 : _GEN_279; // @[TLB.scala 242:54]
  assign _GEN_376 = _T_1077 ? sectored_entries_7_valid_1 : _GEN_280; // @[TLB.scala 242:54]
  assign _GEN_377 = _T_1077 ? sectored_entries_7_valid_2 : _GEN_281; // @[TLB.scala 242:54]
  assign _GEN_378 = _T_1077 ? sectored_entries_7_valid_3 : _GEN_282; // @[TLB.scala 242:54]
  assign _GEN_387 = io_ptw_resp_bits_homogeneous ? special_entry_valid_0 : _GEN_64; // @[TLB.scala 237:68]
  assign _GEN_391 = io_ptw_resp_bits_homogeneous ? _GEN_291 : superpage_entries_0_valid_0; // @[TLB.scala 237:68]
  assign _GEN_395 = io_ptw_resp_bits_homogeneous ? _GEN_295 : superpage_entries_1_valid_0; // @[TLB.scala 237:68]
  assign _GEN_399 = io_ptw_resp_bits_homogeneous ? _GEN_299 : superpage_entries_2_valid_0; // @[TLB.scala 237:68]
  assign _GEN_403 = io_ptw_resp_bits_homogeneous ? _GEN_303 : superpage_entries_3_valid_0; // @[TLB.scala 237:68]
  assign _GEN_405 = io_ptw_resp_bits_homogeneous ? _GEN_305 : sectored_entries_0_valid_0; // @[TLB.scala 237:68]
  assign _GEN_406 = io_ptw_resp_bits_homogeneous ? _GEN_306 : sectored_entries_0_valid_1; // @[TLB.scala 237:68]
  assign _GEN_407 = io_ptw_resp_bits_homogeneous ? _GEN_307 : sectored_entries_0_valid_2; // @[TLB.scala 237:68]
  assign _GEN_408 = io_ptw_resp_bits_homogeneous ? _GEN_308 : sectored_entries_0_valid_3; // @[TLB.scala 237:68]
  assign _GEN_415 = io_ptw_resp_bits_homogeneous ? _GEN_315 : sectored_entries_1_valid_0; // @[TLB.scala 237:68]
  assign _GEN_416 = io_ptw_resp_bits_homogeneous ? _GEN_316 : sectored_entries_1_valid_1; // @[TLB.scala 237:68]
  assign _GEN_417 = io_ptw_resp_bits_homogeneous ? _GEN_317 : sectored_entries_1_valid_2; // @[TLB.scala 237:68]
  assign _GEN_418 = io_ptw_resp_bits_homogeneous ? _GEN_318 : sectored_entries_1_valid_3; // @[TLB.scala 237:68]
  assign _GEN_425 = io_ptw_resp_bits_homogeneous ? _GEN_325 : sectored_entries_2_valid_0; // @[TLB.scala 237:68]
  assign _GEN_426 = io_ptw_resp_bits_homogeneous ? _GEN_326 : sectored_entries_2_valid_1; // @[TLB.scala 237:68]
  assign _GEN_427 = io_ptw_resp_bits_homogeneous ? _GEN_327 : sectored_entries_2_valid_2; // @[TLB.scala 237:68]
  assign _GEN_428 = io_ptw_resp_bits_homogeneous ? _GEN_328 : sectored_entries_2_valid_3; // @[TLB.scala 237:68]
  assign _GEN_435 = io_ptw_resp_bits_homogeneous ? _GEN_335 : sectored_entries_3_valid_0; // @[TLB.scala 237:68]
  assign _GEN_436 = io_ptw_resp_bits_homogeneous ? _GEN_336 : sectored_entries_3_valid_1; // @[TLB.scala 237:68]
  assign _GEN_437 = io_ptw_resp_bits_homogeneous ? _GEN_337 : sectored_entries_3_valid_2; // @[TLB.scala 237:68]
  assign _GEN_438 = io_ptw_resp_bits_homogeneous ? _GEN_338 : sectored_entries_3_valid_3; // @[TLB.scala 237:68]
  assign _GEN_445 = io_ptw_resp_bits_homogeneous ? _GEN_345 : sectored_entries_4_valid_0; // @[TLB.scala 237:68]
  assign _GEN_446 = io_ptw_resp_bits_homogeneous ? _GEN_346 : sectored_entries_4_valid_1; // @[TLB.scala 237:68]
  assign _GEN_447 = io_ptw_resp_bits_homogeneous ? _GEN_347 : sectored_entries_4_valid_2; // @[TLB.scala 237:68]
  assign _GEN_448 = io_ptw_resp_bits_homogeneous ? _GEN_348 : sectored_entries_4_valid_3; // @[TLB.scala 237:68]
  assign _GEN_455 = io_ptw_resp_bits_homogeneous ? _GEN_355 : sectored_entries_5_valid_0; // @[TLB.scala 237:68]
  assign _GEN_456 = io_ptw_resp_bits_homogeneous ? _GEN_356 : sectored_entries_5_valid_1; // @[TLB.scala 237:68]
  assign _GEN_457 = io_ptw_resp_bits_homogeneous ? _GEN_357 : sectored_entries_5_valid_2; // @[TLB.scala 237:68]
  assign _GEN_458 = io_ptw_resp_bits_homogeneous ? _GEN_358 : sectored_entries_5_valid_3; // @[TLB.scala 237:68]
  assign _GEN_465 = io_ptw_resp_bits_homogeneous ? _GEN_365 : sectored_entries_6_valid_0; // @[TLB.scala 237:68]
  assign _GEN_466 = io_ptw_resp_bits_homogeneous ? _GEN_366 : sectored_entries_6_valid_1; // @[TLB.scala 237:68]
  assign _GEN_467 = io_ptw_resp_bits_homogeneous ? _GEN_367 : sectored_entries_6_valid_2; // @[TLB.scala 237:68]
  assign _GEN_468 = io_ptw_resp_bits_homogeneous ? _GEN_368 : sectored_entries_6_valid_3; // @[TLB.scala 237:68]
  assign _GEN_475 = io_ptw_resp_bits_homogeneous ? _GEN_375 : sectored_entries_7_valid_0; // @[TLB.scala 237:68]
  assign _GEN_476 = io_ptw_resp_bits_homogeneous ? _GEN_376 : sectored_entries_7_valid_1; // @[TLB.scala 237:68]
  assign _GEN_477 = io_ptw_resp_bits_homogeneous ? _GEN_377 : sectored_entries_7_valid_2; // @[TLB.scala 237:68]
  assign _GEN_478 = io_ptw_resp_bits_homogeneous ? _GEN_378 : sectored_entries_7_valid_3; // @[TLB.scala 237:68]
  assign _GEN_487 = io_ptw_resp_valid ? _GEN_387 : special_entry_valid_0; // @[TLB.scala 217:20]
  assign _GEN_491 = io_ptw_resp_valid ? _GEN_391 : superpage_entries_0_valid_0; // @[TLB.scala 217:20]
  assign _GEN_495 = io_ptw_resp_valid ? _GEN_395 : superpage_entries_1_valid_0; // @[TLB.scala 217:20]
  assign _GEN_499 = io_ptw_resp_valid ? _GEN_399 : superpage_entries_2_valid_0; // @[TLB.scala 217:20]
  assign _GEN_503 = io_ptw_resp_valid ? _GEN_403 : superpage_entries_3_valid_0; // @[TLB.scala 217:20]
  assign _GEN_505 = io_ptw_resp_valid ? _GEN_405 : sectored_entries_0_valid_0; // @[TLB.scala 217:20]
  assign _GEN_506 = io_ptw_resp_valid ? _GEN_406 : sectored_entries_0_valid_1; // @[TLB.scala 217:20]
  assign _GEN_507 = io_ptw_resp_valid ? _GEN_407 : sectored_entries_0_valid_2; // @[TLB.scala 217:20]
  assign _GEN_508 = io_ptw_resp_valid ? _GEN_408 : sectored_entries_0_valid_3; // @[TLB.scala 217:20]
  assign _GEN_515 = io_ptw_resp_valid ? _GEN_415 : sectored_entries_1_valid_0; // @[TLB.scala 217:20]
  assign _GEN_516 = io_ptw_resp_valid ? _GEN_416 : sectored_entries_1_valid_1; // @[TLB.scala 217:20]
  assign _GEN_517 = io_ptw_resp_valid ? _GEN_417 : sectored_entries_1_valid_2; // @[TLB.scala 217:20]
  assign _GEN_518 = io_ptw_resp_valid ? _GEN_418 : sectored_entries_1_valid_3; // @[TLB.scala 217:20]
  assign _GEN_525 = io_ptw_resp_valid ? _GEN_425 : sectored_entries_2_valid_0; // @[TLB.scala 217:20]
  assign _GEN_526 = io_ptw_resp_valid ? _GEN_426 : sectored_entries_2_valid_1; // @[TLB.scala 217:20]
  assign _GEN_527 = io_ptw_resp_valid ? _GEN_427 : sectored_entries_2_valid_2; // @[TLB.scala 217:20]
  assign _GEN_528 = io_ptw_resp_valid ? _GEN_428 : sectored_entries_2_valid_3; // @[TLB.scala 217:20]
  assign _GEN_535 = io_ptw_resp_valid ? _GEN_435 : sectored_entries_3_valid_0; // @[TLB.scala 217:20]
  assign _GEN_536 = io_ptw_resp_valid ? _GEN_436 : sectored_entries_3_valid_1; // @[TLB.scala 217:20]
  assign _GEN_537 = io_ptw_resp_valid ? _GEN_437 : sectored_entries_3_valid_2; // @[TLB.scala 217:20]
  assign _GEN_538 = io_ptw_resp_valid ? _GEN_438 : sectored_entries_3_valid_3; // @[TLB.scala 217:20]
  assign _GEN_545 = io_ptw_resp_valid ? _GEN_445 : sectored_entries_4_valid_0; // @[TLB.scala 217:20]
  assign _GEN_546 = io_ptw_resp_valid ? _GEN_446 : sectored_entries_4_valid_1; // @[TLB.scala 217:20]
  assign _GEN_547 = io_ptw_resp_valid ? _GEN_447 : sectored_entries_4_valid_2; // @[TLB.scala 217:20]
  assign _GEN_548 = io_ptw_resp_valid ? _GEN_448 : sectored_entries_4_valid_3; // @[TLB.scala 217:20]
  assign _GEN_555 = io_ptw_resp_valid ? _GEN_455 : sectored_entries_5_valid_0; // @[TLB.scala 217:20]
  assign _GEN_556 = io_ptw_resp_valid ? _GEN_456 : sectored_entries_5_valid_1; // @[TLB.scala 217:20]
  assign _GEN_557 = io_ptw_resp_valid ? _GEN_457 : sectored_entries_5_valid_2; // @[TLB.scala 217:20]
  assign _GEN_558 = io_ptw_resp_valid ? _GEN_458 : sectored_entries_5_valid_3; // @[TLB.scala 217:20]
  assign _GEN_565 = io_ptw_resp_valid ? _GEN_465 : sectored_entries_6_valid_0; // @[TLB.scala 217:20]
  assign _GEN_566 = io_ptw_resp_valid ? _GEN_466 : sectored_entries_6_valid_1; // @[TLB.scala 217:20]
  assign _GEN_567 = io_ptw_resp_valid ? _GEN_467 : sectored_entries_6_valid_2; // @[TLB.scala 217:20]
  assign _GEN_568 = io_ptw_resp_valid ? _GEN_468 : sectored_entries_6_valid_3; // @[TLB.scala 217:20]
  assign _GEN_575 = io_ptw_resp_valid ? _GEN_475 : sectored_entries_7_valid_0; // @[TLB.scala 217:20]
  assign _GEN_576 = io_ptw_resp_valid ? _GEN_476 : sectored_entries_7_valid_1; // @[TLB.scala 217:20]
  assign _GEN_577 = io_ptw_resp_valid ? _GEN_477 : sectored_entries_7_valid_2; // @[TLB.scala 217:20]
  assign _GEN_578 = io_ptw_resp_valid ? _GEN_478 : sectored_entries_7_valid_3; // @[TLB.scala 217:20]
  assign _T_1761 = {OptimizationBarrier_19_io_y_ae,OptimizationBarrier_18_io_y_ae,OptimizationBarrier_17_io_y_ae,OptimizationBarrier_16_io_y_ae,OptimizationBarrier_15_io_y_ae,OptimizationBarrier_14_io_y_ae}; // @[Cat.scala 29:58]
  assign ptw_ae_array = {1'h0,OptimizationBarrier_26_io_y_ae,OptimizationBarrier_25_io_y_ae,OptimizationBarrier_24_io_y_ae,OptimizationBarrier_23_io_y_ae,OptimizationBarrier_22_io_y_ae,OptimizationBarrier_21_io_y_ae,OptimizationBarrier_20_io_y_ae,_T_1761}; // @[Cat.scala 29:58]
  assign _T_1770 = ~priv_s | io_ptw_status_sum; // @[TLB.scala 261:32]
  assign _T_1775 = {OptimizationBarrier_19_io_y_u,OptimizationBarrier_18_io_y_u,OptimizationBarrier_17_io_y_u,OptimizationBarrier_16_io_y_u,OptimizationBarrier_15_io_y_u,OptimizationBarrier_14_io_y_u}; // @[Cat.scala 29:58]
  assign _T_1782 = {OptimizationBarrier_26_io_y_u,OptimizationBarrier_25_io_y_u,OptimizationBarrier_24_io_y_u,OptimizationBarrier_23_io_y_u,OptimizationBarrier_22_io_y_u,OptimizationBarrier_21_io_y_u,OptimizationBarrier_20_io_y_u,_T_1775}; // @[Cat.scala 29:58]
  assign _T_1783 = _T_1770 ? _T_1782 : 13'h0; // @[TLB.scala 261:23]
  assign _T_1797 = priv_s ? ~_T_1782 : 13'h0; // @[TLB.scala 261:89]
  assign priv_rw_ok = _T_1783 | _T_1797; // @[TLB.scala 261:84]
  assign _T_1827 = {OptimizationBarrier_19_io_y_sr,OptimizationBarrier_18_io_y_sr,OptimizationBarrier_17_io_y_sr,OptimizationBarrier_16_io_y_sr,OptimizationBarrier_15_io_y_sr,OptimizationBarrier_14_io_y_sr}; // @[Cat.scala 29:58]
  assign _T_1834 = {OptimizationBarrier_26_io_y_sr,OptimizationBarrier_25_io_y_sr,OptimizationBarrier_24_io_y_sr,OptimizationBarrier_23_io_y_sr,OptimizationBarrier_22_io_y_sr,OptimizationBarrier_21_io_y_sr,OptimizationBarrier_20_io_y_sr,_T_1827}; // @[Cat.scala 29:58]
  assign _T_1839 = {OptimizationBarrier_19_io_y_sx,OptimizationBarrier_18_io_y_sx,OptimizationBarrier_17_io_y_sx,OptimizationBarrier_16_io_y_sx,OptimizationBarrier_15_io_y_sx,OptimizationBarrier_14_io_y_sx}; // @[Cat.scala 29:58]
  assign _T_1846 = {OptimizationBarrier_26_io_y_sx,OptimizationBarrier_25_io_y_sx,OptimizationBarrier_24_io_y_sx,OptimizationBarrier_23_io_y_sx,OptimizationBarrier_22_io_y_sx,OptimizationBarrier_21_io_y_sx,OptimizationBarrier_20_io_y_sx,_T_1839}; // @[Cat.scala 29:58]
  assign _T_1847 = io_ptw_status_mxr ? _T_1846 : 13'h0; // @[TLB.scala 263:73]
  assign _T_1848 = _T_1834 | _T_1847; // @[TLB.scala 263:68]
  assign _T_1849 = priv_rw_ok & _T_1848; // @[TLB.scala 263:40]
  assign r_array = {1'h1,_T_1849}; // @[Cat.scala 29:58]
  assign _T_1854 = {OptimizationBarrier_19_io_y_sw,OptimizationBarrier_18_io_y_sw,OptimizationBarrier_17_io_y_sw,OptimizationBarrier_16_io_y_sw,OptimizationBarrier_15_io_y_sw,OptimizationBarrier_14_io_y_sw}; // @[Cat.scala 29:58]
  assign _T_1861 = {OptimizationBarrier_26_io_y_sw,OptimizationBarrier_25_io_y_sw,OptimizationBarrier_24_io_y_sw,OptimizationBarrier_23_io_y_sw,OptimizationBarrier_22_io_y_sw,OptimizationBarrier_21_io_y_sw,OptimizationBarrier_20_io_y_sw,_T_1854}; // @[Cat.scala 29:58]
  assign _T_1862 = priv_rw_ok & _T_1861; // @[TLB.scala 264:40]
  assign w_array = {1'h1,_T_1862}; // @[Cat.scala 29:58]
  assign _T_1877 = prot_r ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_1882 = {OptimizationBarrier_32_io_y_pr,OptimizationBarrier_31_io_y_pr,OptimizationBarrier_30_io_y_pr,OptimizationBarrier_29_io_y_pr,OptimizationBarrier_28_io_y_pr,OptimizationBarrier_27_io_y_pr}; // @[Cat.scala 29:58]
  assign _T_1889 = {_T_1877,OptimizationBarrier_38_io_y_pr,OptimizationBarrier_37_io_y_pr,OptimizationBarrier_36_io_y_pr,OptimizationBarrier_35_io_y_pr,OptimizationBarrier_34_io_y_pr,OptimizationBarrier_33_io_y_pr,_T_1882}; // @[Cat.scala 29:58]
  assign pr_array = _T_1889 & ~ptw_ae_array; // @[TLB.scala 266:87]
  assign _T_1892 = prot_w ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_1897 = {OptimizationBarrier_32_io_y_pw,OptimizationBarrier_31_io_y_pw,OptimizationBarrier_30_io_y_pw,OptimizationBarrier_29_io_y_pw,OptimizationBarrier_28_io_y_pw,OptimizationBarrier_27_io_y_pw}; // @[Cat.scala 29:58]
  assign _T_1904 = {_T_1892,OptimizationBarrier_38_io_y_pw,OptimizationBarrier_37_io_y_pw,OptimizationBarrier_36_io_y_pw,OptimizationBarrier_35_io_y_pw,OptimizationBarrier_34_io_y_pw,OptimizationBarrier_33_io_y_pw,_T_1897}; // @[Cat.scala 29:58]
  assign pw_array = _T_1904 & ~ptw_ae_array; // @[TLB.scala 267:87]
  assign _T_1922 = prot_eff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_1927 = {OptimizationBarrier_32_io_y_eff,OptimizationBarrier_31_io_y_eff,OptimizationBarrier_30_io_y_eff,OptimizationBarrier_29_io_y_eff,OptimizationBarrier_28_io_y_eff,OptimizationBarrier_27_io_y_eff}; // @[Cat.scala 29:58]
  assign eff_array = {_T_1922,OptimizationBarrier_38_io_y_eff,OptimizationBarrier_37_io_y_eff,OptimizationBarrier_36_io_y_eff,OptimizationBarrier_35_io_y_eff,OptimizationBarrier_34_io_y_eff,OptimizationBarrier_33_io_y_eff,_T_1927}; // @[Cat.scala 29:58]
  assign _T_1935 = cacheable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_1940 = {OptimizationBarrier_32_io_y_c,OptimizationBarrier_31_io_y_c,OptimizationBarrier_30_io_y_c,OptimizationBarrier_29_io_y_c,OptimizationBarrier_28_io_y_c,OptimizationBarrier_27_io_y_c}; // @[Cat.scala 29:58]
  assign c_array = {_T_1935,OptimizationBarrier_38_io_y_c,OptimizationBarrier_37_io_y_c,OptimizationBarrier_36_io_y_c,OptimizationBarrier_35_io_y_c,OptimizationBarrier_34_io_y_c,OptimizationBarrier_33_io_y_c,_T_1940}; // @[Cat.scala 29:58]
  assign _T_1948 = _T_239 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_1953 = {OptimizationBarrier_32_io_y_ppp,OptimizationBarrier_31_io_y_ppp,OptimizationBarrier_30_io_y_ppp,OptimizationBarrier_29_io_y_ppp,OptimizationBarrier_28_io_y_ppp,OptimizationBarrier_27_io_y_ppp}; // @[Cat.scala 29:58]
  assign ppp_array = {_T_1948,OptimizationBarrier_38_io_y_ppp,OptimizationBarrier_37_io_y_ppp,OptimizationBarrier_36_io_y_ppp,OptimizationBarrier_35_io_y_ppp,OptimizationBarrier_34_io_y_ppp,OptimizationBarrier_33_io_y_ppp,_T_1953}; // @[Cat.scala 29:58]
  assign _T_1961 = prot_al ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_1966 = {OptimizationBarrier_32_io_y_paa,OptimizationBarrier_31_io_y_paa,OptimizationBarrier_30_io_y_paa,OptimizationBarrier_29_io_y_paa,OptimizationBarrier_28_io_y_paa,OptimizationBarrier_27_io_y_paa}; // @[Cat.scala 29:58]
  assign paa_array = {_T_1961,OptimizationBarrier_38_io_y_paa,OptimizationBarrier_37_io_y_paa,OptimizationBarrier_36_io_y_paa,OptimizationBarrier_35_io_y_paa,OptimizationBarrier_34_io_y_paa,OptimizationBarrier_33_io_y_paa,_T_1966}; // @[Cat.scala 29:58]
  assign _T_1979 = {OptimizationBarrier_32_io_y_pal,OptimizationBarrier_31_io_y_pal,OptimizationBarrier_30_io_y_pal,OptimizationBarrier_29_io_y_pal,OptimizationBarrier_28_io_y_pal,OptimizationBarrier_27_io_y_pal}; // @[Cat.scala 29:58]
  assign pal_array = {_T_1961,OptimizationBarrier_38_io_y_pal,OptimizationBarrier_37_io_y_pal,OptimizationBarrier_36_io_y_pal,OptimizationBarrier_35_io_y_pal,OptimizationBarrier_34_io_y_pal,OptimizationBarrier_33_io_y_pal,_T_1979}; // @[Cat.scala 29:58]
  assign ppp_array_if_cached = ppp_array | c_array; // @[TLB.scala 274:39]
  assign paa_array_if_cached = paa_array | c_array; // @[TLB.scala 275:39]
  assign pal_array_if_cached = pal_array | c_array; // @[TLB.scala 276:39]
  assign _T_2001 = 4'h1 << io_req_bits_size; // @[OneHot.scala 58:35]
  assign _T_2003 = _T_2001 - 4'h1; // @[TLB.scala 279:69]
  assign _GEN_1027 = {{36'd0}, _T_2003}; // @[TLB.scala 279:39]
  assign _T_2004 = io_req_bits_vaddr & _GEN_1027; // @[TLB.scala 279:39]
  assign misaligned = |_T_2004; // @[TLB.scala 279:75]
  assign _T_2005 = io_req_bits_vaddr & 40'hc000000000; // @[TLB.scala 285:43]
  assign _T_2007 = _T_2005 == 40'h0; // @[TLB.scala 286:61]
  assign _T_2008 = _T_2005 == 40'hc000000000; // @[TLB.scala 286:82]
  assign _T_2009 = _T_2007 | _T_2008; // @[TLB.scala 286:67]
  assign bad_va = vm_enabled & ~_T_2009; // @[TLB.scala 280:117]
  assign _T_2012 = io_req_bits_cmd == 5'h6; // @[package.scala 15:47]
  assign _T_2013 = io_req_bits_cmd == 5'h7; // @[package.scala 15:47]
  assign cmd_lrsc = _T_2012 | _T_2013; // @[package.scala 64:59]
  assign _T_2015 = io_req_bits_cmd == 5'h4; // @[package.scala 15:47]
  assign _T_2016 = io_req_bits_cmd == 5'h9; // @[package.scala 15:47]
  assign _T_2017 = io_req_bits_cmd == 5'ha; // @[package.scala 15:47]
  assign _T_2018 = io_req_bits_cmd == 5'hb; // @[package.scala 15:47]
  assign _T_2019 = _T_2015 | _T_2016; // @[package.scala 64:59]
  assign _T_2020 = _T_2019 | _T_2017; // @[package.scala 64:59]
  assign cmd_amo_logical = _T_2020 | _T_2018; // @[package.scala 64:59]
  assign _T_2022 = io_req_bits_cmd == 5'h8; // @[package.scala 15:47]
  assign _T_2023 = io_req_bits_cmd == 5'hc; // @[package.scala 15:47]
  assign _T_2024 = io_req_bits_cmd == 5'hd; // @[package.scala 15:47]
  assign _T_2025 = io_req_bits_cmd == 5'he; // @[package.scala 15:47]
  assign _T_2026 = io_req_bits_cmd == 5'hf; // @[package.scala 15:47]
  assign _T_2027 = _T_2022 | _T_2023; // @[package.scala 64:59]
  assign _T_2028 = _T_2027 | _T_2024; // @[package.scala 64:59]
  assign _T_2029 = _T_2028 | _T_2025; // @[package.scala 64:59]
  assign cmd_amo_arithmetic = _T_2029 | _T_2026; // @[package.scala 64:59]
  assign cmd_put_partial = io_req_bits_cmd == 5'h11; // @[TLB.scala 293:41]
  assign _T_2031 = io_req_bits_cmd == 5'h0; // @[Consts.scala 82:31]
  assign _T_2033 = _T_2031 | _T_2012; // @[Consts.scala 82:41]
  assign _T_2035 = _T_2033 | _T_2013; // @[Consts.scala 82:58]
  assign _T_2052 = cmd_amo_logical | cmd_amo_arithmetic; // @[Consts.scala 80:44]
  assign cmd_read = _T_2035 | _T_2052; // @[Consts.scala 82:75]
  assign _T_2053 = io_req_bits_cmd == 5'h1; // @[Consts.scala 83:32]
  assign _T_2055 = _T_2053 | cmd_put_partial; // @[Consts.scala 83:42]
  assign _T_2057 = _T_2055 | _T_2013; // @[Consts.scala 83:59]
  assign cmd_write = _T_2057 | _T_2052; // @[Consts.scala 83:76]
  assign _T_2075 = io_req_bits_cmd == 5'h5; // @[package.scala 15:47]
  assign _T_2076 = io_req_bits_cmd == 5'h17; // @[package.scala 15:47]
  assign _T_2077 = _T_2075 | _T_2076; // @[package.scala 64:59]
  assign cmd_write_perms = cmd_write | _T_2077; // @[TLB.scala 296:35]
  assign _T_2078 = misaligned ? eff_array : 14'h0; // @[TLB.scala 301:8]
  assign _T_2080 = cmd_lrsc ? ~c_array : 14'h0; // @[TLB.scala 302:8]
  assign ae_array = _T_2078 | _T_2080; // @[TLB.scala 301:37]
  assign _T_2082 = ae_array | ~pr_array; // @[TLB.scala 303:44]
  assign ae_ld_array = cmd_read ? _T_2082 : 14'h0; // @[TLB.scala 303:24]
  assign _T_2084 = ae_array | ~pw_array; // @[TLB.scala 305:35]
  assign _T_2085 = cmd_write_perms ? _T_2084 : 14'h0; // @[TLB.scala 305:8]
  assign _T_2087 = cmd_put_partial ? ~ppp_array_if_cached : 14'h0; // @[TLB.scala 306:8]
  assign _T_2088 = _T_2085 | _T_2087; // @[TLB.scala 305:53]
  assign _T_2090 = cmd_amo_logical ? ~pal_array_if_cached : 14'h0; // @[TLB.scala 307:8]
  assign _T_2091 = _T_2088 | _T_2090; // @[TLB.scala 306:53]
  assign _T_2093 = cmd_amo_arithmetic ? ~paa_array_if_cached : 14'h0; // @[TLB.scala 308:8]
  assign ae_st_array = _T_2091 | _T_2093; // @[TLB.scala 307:53]
  assign _T_2104 = misaligned & cmd_read; // @[TLB.scala 314:36]
  assign ma_ld_array = _T_2104 ? ~eff_array : 14'h0; // @[TLB.scala 314:24]
  assign _T_2106 = misaligned & cmd_write; // @[TLB.scala 315:36]
  assign ma_st_array = _T_2106 ? ~eff_array : 14'h0; // @[TLB.scala 315:24]
  assign _T_2108 = r_array | ptw_ae_array; // @[TLB.scala 316:45]
  assign pf_ld_array = cmd_read ? ~_T_2108 : 14'h0; // @[TLB.scala 316:24]
  assign _T_2110 = w_array | ptw_ae_array; // @[TLB.scala 317:52]
  assign pf_st_array = cmd_write_perms ? ~_T_2110 : 14'h0; // @[TLB.scala 317:24]
  assign tlb_hit = |real_hits; // @[TLB.scala 320:27]
  assign _T_2114 = vm_enabled & ~bad_va; // @[TLB.scala 321:29]
  assign tlb_miss = _T_2114 & ~tlb_hit; // @[TLB.scala 321:40]
  assign _T_2118 = io_req_valid & vm_enabled; // @[TLB.scala 325:22]
  assign _T_2119 = sector_hits_0 | sector_hits_1; // @[package.scala 64:59]
  assign _T_2120 = _T_2119 | sector_hits_2; // @[package.scala 64:59]
  assign _T_2121 = _T_2120 | sector_hits_3; // @[package.scala 64:59]
  assign _T_2122 = _T_2121 | sector_hits_4; // @[package.scala 64:59]
  assign _T_2123 = _T_2122 | sector_hits_5; // @[package.scala 64:59]
  assign _T_2124 = _T_2123 | sector_hits_6; // @[package.scala 64:59]
  assign _T_2125 = _T_2124 | sector_hits_7; // @[package.scala 64:59]
  assign _T_2132 = {sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0}; // @[Cat.scala 29:58]
  assign _T_2135 = |_T_2132[7:4]; // @[OneHot.scala 32:14]
  assign _T_2136 = _T_2132[7:4] | _T_2132[3:0]; // @[OneHot.scala 32:28]
  assign _T_2139 = |_T_2136[3:2]; // @[OneHot.scala 32:14]
  assign _T_2140 = _T_2136[3:2] | _T_2136[1:0]; // @[OneHot.scala 32:28]
  assign _T_2143 = {_T_2135,_T_2139,_T_2140[1]}; // @[Cat.scala 29:58]
  assign _T_2157 = _T_2143[1] ? ~_T_2143[0] : _T_2116[4]; // @[Replacement.scala 193:16]
  assign _T_2161 = _T_2143[1] ? _T_2116[3] : ~_T_2143[0]; // @[Replacement.scala 196:16]
  assign _T_2163 = {~_T_2143[1],_T_2157,_T_2161}; // @[Cat.scala 29:58]
  assign _T_2164 = _T_2143[2] ? _T_2163 : _T_2116[5:3]; // @[Replacement.scala 193:16]
  assign _T_2173 = _T_2143[1] ? ~_T_2143[0] : _T_2116[1]; // @[Replacement.scala 193:16]
  assign _T_2177 = _T_2143[1] ? _T_2116[0] : ~_T_2143[0]; // @[Replacement.scala 196:16]
  assign _T_2179 = {~_T_2143[1],_T_2173,_T_2177}; // @[Cat.scala 29:58]
  assign _T_2180 = _T_2143[2] ? _T_2116[2:0] : _T_2179; // @[Replacement.scala 196:16]
  assign _T_2182 = {~_T_2143[2],_T_2164,_T_2180}; // @[Cat.scala 29:58]
  assign _T_2183 = superpage_hits_0 | superpage_hits_1; // @[package.scala 64:59]
  assign _T_2184 = _T_2183 | superpage_hits_2; // @[package.scala 64:59]
  assign _T_2185 = _T_2184 | superpage_hits_3; // @[package.scala 64:59]
  assign _T_2188 = {superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; // @[Cat.scala 29:58]
  assign _T_2191 = |_T_2188[3:2]; // @[OneHot.scala 32:14]
  assign _T_2192 = _T_2188[3:2] | _T_2188[1:0]; // @[OneHot.scala 32:28]
  assign _T_2194 = {_T_2191,_T_2192[1]}; // @[Cat.scala 29:58]
  assign _T_2203 = _T_2194[1] ? ~_T_2194[0] : _T_2117[1]; // @[Replacement.scala 193:16]
  assign _T_2207 = _T_2194[1] ? _T_2117[0] : ~_T_2194[0]; // @[Replacement.scala 196:16]
  assign _T_2209 = {~_T_2194[1],_T_2203,_T_2207}; // @[Cat.scala 29:58]
  assign _T_2219 = real_hits[1] | real_hits[2]; // @[Misc.scala 182:16]
  assign _T_2221 = real_hits[1] & real_hits[2]; // @[Misc.scala 182:61]
  assign _T_2223 = real_hits[0] | _T_2219; // @[Misc.scala 182:16]
  assign _T_2225 = real_hits[0] & _T_2219; // @[Misc.scala 182:61]
  assign _T_2226 = _T_2221 | _T_2225; // @[Misc.scala 182:49]
  assign _T_2235 = real_hits[4] | real_hits[5]; // @[Misc.scala 182:16]
  assign _T_2237 = real_hits[4] & real_hits[5]; // @[Misc.scala 182:61]
  assign _T_2239 = real_hits[3] | _T_2235; // @[Misc.scala 182:16]
  assign _T_2241 = real_hits[3] & _T_2235; // @[Misc.scala 182:61]
  assign _T_2242 = _T_2237 | _T_2241; // @[Misc.scala 182:49]
  assign _T_2243 = _T_2223 | _T_2239; // @[Misc.scala 182:16]
  assign _T_2244 = _T_2226 | _T_2242; // @[Misc.scala 182:37]
  assign _T_2245 = _T_2223 & _T_2239; // @[Misc.scala 182:61]
  assign _T_2246 = _T_2244 | _T_2245; // @[Misc.scala 182:49]
  assign _T_2256 = real_hits[7] | real_hits[8]; // @[Misc.scala 182:16]
  assign _T_2258 = real_hits[7] & real_hits[8]; // @[Misc.scala 182:61]
  assign _T_2260 = real_hits[6] | _T_2256; // @[Misc.scala 182:16]
  assign _T_2262 = real_hits[6] & _T_2256; // @[Misc.scala 182:61]
  assign _T_2263 = _T_2258 | _T_2262; // @[Misc.scala 182:49]
  assign _T_2270 = real_hits[9] | real_hits[10]; // @[Misc.scala 182:16]
  assign _T_2272 = real_hits[9] & real_hits[10]; // @[Misc.scala 182:61]
  assign _T_2279 = real_hits[11] | real_hits[12]; // @[Misc.scala 182:16]
  assign _T_2281 = real_hits[11] & real_hits[12]; // @[Misc.scala 182:61]
  assign _T_2283 = _T_2270 | _T_2279; // @[Misc.scala 182:16]
  assign _T_2284 = _T_2272 | _T_2281; // @[Misc.scala 182:37]
  assign _T_2285 = _T_2270 & _T_2279; // @[Misc.scala 182:61]
  assign _T_2286 = _T_2284 | _T_2285; // @[Misc.scala 182:49]
  assign _T_2287 = _T_2260 | _T_2283; // @[Misc.scala 182:16]
  assign _T_2288 = _T_2263 | _T_2286; // @[Misc.scala 182:37]
  assign _T_2289 = _T_2260 & _T_2283; // @[Misc.scala 182:61]
  assign _T_2290 = _T_2288 | _T_2289; // @[Misc.scala 182:49]
  assign _T_2292 = _T_2246 | _T_2290; // @[Misc.scala 182:37]
  assign _T_2293 = _T_2243 & _T_2287; // @[Misc.scala 182:61]
  assign multipleHits = _T_2292 | _T_2293; // @[Misc.scala 182:49]
  assign _T_2295 = bad_va & cmd_read; // @[TLB.scala 338:28]
  assign _T_2296 = pf_ld_array & hits; // @[TLB.scala 338:57]
  assign _T_2297 = |_T_2296; // @[TLB.scala 338:65]
  assign _T_2299 = bad_va & cmd_write_perms; // @[TLB.scala 339:28]
  assign _T_2300 = pf_st_array & hits; // @[TLB.scala 339:64]
  assign _T_2301 = |_T_2300; // @[TLB.scala 339:72]
  assign _T_2306 = ae_ld_array & hits; // @[TLB.scala 341:33]
  assign _T_2308 = ae_st_array & hits; // @[TLB.scala 342:33]
  assign _T_2313 = ma_ld_array & hits; // @[TLB.scala 344:33]
  assign _T_2315 = ma_st_array & hits; // @[TLB.scala 345:33]
  assign _T_2317 = c_array & hits; // @[TLB.scala 347:33]
  assign _T_2324 = io_ptw_resp_valid | tlb_miss; // @[TLB.scala 350:29]
  assign _T_2330 = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37]
  assign _T_2331 = _T_2330 & tlb_miss; // @[TLB.scala 359:25]
  assign _T_2337 = _T_2117[2] ? _T_2117[1] : _T_2117[0]; // @[Replacement.scala 240:16]
  assign _T_2338 = {_T_2117[2],_T_2337}; // @[Cat.scala 29:58]
  assign _T_2341 = {superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[Cat.scala 29:58]
  assign _T_2342 = &_T_2341; // @[TLB.scala 407:16]
  assign _T_2344 = ~_T_2341[0]; // @[OneHot.scala 47:40]
  assign _T_2345 = ~_T_2341[1]; // @[OneHot.scala 47:40]
  assign _T_2346 = ~_T_2341[2]; // @[OneHot.scala 47:40]
  assign _T_2360 = _T_2116[5] ? _T_2116[4] : _T_2116[3]; // @[Replacement.scala 240:16]
  assign _T_2361 = {_T_2116[5],_T_2360}; // @[Cat.scala 29:58]
  assign _T_2367 = _T_2116[2] ? _T_2116[1] : _T_2116[0]; // @[Replacement.scala 240:16]
  assign _T_2368 = {_T_2116[2],_T_2367}; // @[Cat.scala 29:58]
  assign _T_2369 = _T_2116[6] ? _T_2361 : _T_2368; // @[Replacement.scala 240:16]
  assign _T_2370 = {_T_2116[6],_T_2369}; // @[Cat.scala 29:58]
  assign _T_2401 = {_T_461,_T_455,_T_449,_T_443,_T_437,_T_431,_T_425,_T_419}; // @[Cat.scala 29:58]
  assign _T_2402 = &_T_2401; // @[TLB.scala 407:16]
  assign _T_2404 = ~_T_2401[0]; // @[OneHot.scala 47:40]
  assign _T_2405 = ~_T_2401[1]; // @[OneHot.scala 47:40]
  assign _T_2406 = ~_T_2401[2]; // @[OneHot.scala 47:40]
  assign _T_2407 = ~_T_2401[3]; // @[OneHot.scala 47:40]
  assign _T_2408 = ~_T_2401[4]; // @[OneHot.scala 47:40]
  assign _T_2409 = ~_T_2401[5]; // @[OneHot.scala 47:40]
  assign _T_2410 = ~_T_2401[6]; // @[OneHot.scala 47:40]
  assign _T_2447 = state == 2'h2; // @[TLB.scala 373:17]
  assign _T_2448 = _T_2447 & io_sfence_valid; // @[TLB.scala 373:28]
  assign _T_2451 = io_sfence_bits_addr[38:12] == vpn; // @[TLB.scala 381:72]
  assign _T_2452 = ~io_sfence_bits_rs1 | _T_2451; // @[TLB.scala 381:34]
  assign _T_2454 = _T_2452 | reset; // @[TLB.scala 381:13]
  assign _T_2462 = _T_420[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_681 = sectored_entries_0_data_0[13] ? _GEN_505 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_682 = sectored_entries_0_data_1[13] ? _GEN_506 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_683 = sectored_entries_0_data_2[13] ? _GEN_507 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_684 = sectored_entries_0_data_3[13] ? _GEN_508 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_685 = io_sfence_bits_rs2 & _GEN_681; // @[TLB.scala 384:40]
  assign _GEN_686 = io_sfence_bits_rs2 & _GEN_682; // @[TLB.scala 384:40]
  assign _GEN_687 = io_sfence_bits_rs2 & _GEN_683; // @[TLB.scala 384:40]
  assign _GEN_688 = io_sfence_bits_rs2 & _GEN_684; // @[TLB.scala 384:40]
  assign _T_2617 = _T_426[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_709 = sectored_entries_1_data_0[13] ? _GEN_515 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_710 = sectored_entries_1_data_1[13] ? _GEN_516 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_711 = sectored_entries_1_data_2[13] ? _GEN_517 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_712 = sectored_entries_1_data_3[13] ? _GEN_518 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_713 = io_sfence_bits_rs2 & _GEN_709; // @[TLB.scala 384:40]
  assign _GEN_714 = io_sfence_bits_rs2 & _GEN_710; // @[TLB.scala 384:40]
  assign _GEN_715 = io_sfence_bits_rs2 & _GEN_711; // @[TLB.scala 384:40]
  assign _GEN_716 = io_sfence_bits_rs2 & _GEN_712; // @[TLB.scala 384:40]
  assign _T_2772 = _T_432[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_737 = sectored_entries_2_data_0[13] ? _GEN_525 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_738 = sectored_entries_2_data_1[13] ? _GEN_526 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_739 = sectored_entries_2_data_2[13] ? _GEN_527 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_740 = sectored_entries_2_data_3[13] ? _GEN_528 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_741 = io_sfence_bits_rs2 & _GEN_737; // @[TLB.scala 384:40]
  assign _GEN_742 = io_sfence_bits_rs2 & _GEN_738; // @[TLB.scala 384:40]
  assign _GEN_743 = io_sfence_bits_rs2 & _GEN_739; // @[TLB.scala 384:40]
  assign _GEN_744 = io_sfence_bits_rs2 & _GEN_740; // @[TLB.scala 384:40]
  assign _T_2927 = _T_438[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_765 = sectored_entries_3_data_0[13] ? _GEN_535 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_766 = sectored_entries_3_data_1[13] ? _GEN_536 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_767 = sectored_entries_3_data_2[13] ? _GEN_537 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_768 = sectored_entries_3_data_3[13] ? _GEN_538 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_769 = io_sfence_bits_rs2 & _GEN_765; // @[TLB.scala 384:40]
  assign _GEN_770 = io_sfence_bits_rs2 & _GEN_766; // @[TLB.scala 384:40]
  assign _GEN_771 = io_sfence_bits_rs2 & _GEN_767; // @[TLB.scala 384:40]
  assign _GEN_772 = io_sfence_bits_rs2 & _GEN_768; // @[TLB.scala 384:40]
  assign _T_3082 = _T_444[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_793 = sectored_entries_4_data_0[13] ? _GEN_545 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_794 = sectored_entries_4_data_1[13] ? _GEN_546 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_795 = sectored_entries_4_data_2[13] ? _GEN_547 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_796 = sectored_entries_4_data_3[13] ? _GEN_548 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_797 = io_sfence_bits_rs2 & _GEN_793; // @[TLB.scala 384:40]
  assign _GEN_798 = io_sfence_bits_rs2 & _GEN_794; // @[TLB.scala 384:40]
  assign _GEN_799 = io_sfence_bits_rs2 & _GEN_795; // @[TLB.scala 384:40]
  assign _GEN_800 = io_sfence_bits_rs2 & _GEN_796; // @[TLB.scala 384:40]
  assign _T_3237 = _T_450[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_821 = sectored_entries_5_data_0[13] ? _GEN_555 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_822 = sectored_entries_5_data_1[13] ? _GEN_556 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_823 = sectored_entries_5_data_2[13] ? _GEN_557 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_824 = sectored_entries_5_data_3[13] ? _GEN_558 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_825 = io_sfence_bits_rs2 & _GEN_821; // @[TLB.scala 384:40]
  assign _GEN_826 = io_sfence_bits_rs2 & _GEN_822; // @[TLB.scala 384:40]
  assign _GEN_827 = io_sfence_bits_rs2 & _GEN_823; // @[TLB.scala 384:40]
  assign _GEN_828 = io_sfence_bits_rs2 & _GEN_824; // @[TLB.scala 384:40]
  assign _T_3392 = _T_456[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_849 = sectored_entries_6_data_0[13] ? _GEN_565 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_850 = sectored_entries_6_data_1[13] ? _GEN_566 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_851 = sectored_entries_6_data_2[13] ? _GEN_567 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_852 = sectored_entries_6_data_3[13] ? _GEN_568 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_853 = io_sfence_bits_rs2 & _GEN_849; // @[TLB.scala 384:40]
  assign _GEN_854 = io_sfence_bits_rs2 & _GEN_850; // @[TLB.scala 384:40]
  assign _GEN_855 = io_sfence_bits_rs2 & _GEN_851; // @[TLB.scala 384:40]
  assign _GEN_856 = io_sfence_bits_rs2 & _GEN_852; // @[TLB.scala 384:40]
  assign _T_3547 = _T_462[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_877 = sectored_entries_7_data_0[13] ? _GEN_575 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_878 = sectored_entries_7_data_1[13] ? _GEN_576 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_879 = sectored_entries_7_data_2[13] ? _GEN_577 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_880 = sectored_entries_7_data_3[13] ? _GEN_578 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_881 = io_sfence_bits_rs2 & _GEN_877; // @[TLB.scala 384:40]
  assign _GEN_882 = io_sfence_bits_rs2 & _GEN_878; // @[TLB.scala 384:40]
  assign _GEN_883 = io_sfence_bits_rs2 & _GEN_879; // @[TLB.scala 384:40]
  assign _GEN_884 = io_sfence_bits_rs2 & _GEN_880; // @[TLB.scala 384:40]
  assign _GEN_890 = superpage_entries_0_data_0[13] ? _GEN_491 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_891 = io_sfence_bits_rs2 & _GEN_890; // @[TLB.scala 384:40]
  assign _GEN_894 = superpage_entries_1_data_0[13] ? _GEN_495 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_895 = io_sfence_bits_rs2 & _GEN_894; // @[TLB.scala 384:40]
  assign _GEN_898 = superpage_entries_2_data_0[13] ? _GEN_499 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_899 = io_sfence_bits_rs2 & _GEN_898; // @[TLB.scala 384:40]
  assign _GEN_902 = superpage_entries_3_data_0[13] ? _GEN_503 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_903 = io_sfence_bits_rs2 & _GEN_902; // @[TLB.scala 384:40]
  assign _GEN_906 = special_entry_data_0[13] ? _GEN_487 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_907 = io_sfence_bits_rs2 & _GEN_906; // @[TLB.scala 384:40]
  assign _T_3897 = multipleHits | reset; // @[TLB.scala 388:24]
  assign io_req_ready = state == 2'h0; // @[TLB.scala 337:16]
  assign io_resp_miss = _T_2324 | multipleHits; // @[TLB.scala 350:16]
  assign io_resp_paddr = {ppn,io_req_bits_vaddr[11:0]}; // @[TLB.scala 351:17]
  assign io_resp_pf_ld = _T_2295 | _T_2297; // @[TLB.scala 338:17]
  assign io_resp_pf_st = _T_2299 | _T_2301; // @[TLB.scala 339:17]
  assign io_resp_ae_ld = |_T_2306; // @[TLB.scala 341:17]
  assign io_resp_ae_st = |_T_2308; // @[TLB.scala 342:17]
  assign io_resp_ma_ld = |_T_2313; // @[TLB.scala 344:17]
  assign io_resp_ma_st = |_T_2315; // @[TLB.scala 345:17]
  assign io_resp_cacheable = |_T_2317; // @[TLB.scala 347:21]
  assign io_ptw_req_valid = state == 2'h1; // @[TLB.scala 353:20]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[TLB.scala 355:29]
  assign OptimizationBarrier_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_u = special_entry_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_ae = special_entry_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_sw = special_entry_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_sx = special_entry_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_sr = special_entry_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_pw = special_entry_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_px = special_entry_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_pr = special_entry_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_ppp = special_entry_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_pal = special_entry_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_paa = special_entry_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_eff = special_entry_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_c = special_entry_data_0[1]; // @[package.scala 244:18]
  assign pmp_io_prv = mpu_priv[1:0]; // @[TLB.scala 194:14]
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask; // @[TLB.scala 193:14]
  assign pmp_io_addr = mpu_physaddr[31:0]; // @[TLB.scala 191:15]
  assign pmp_io_size = io_req_bits_size; // @[TLB.scala 192:15]
  assign OptimizationBarrier_1_io_x_ppn = _GEN_35[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_u = _GEN_35[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_ae = _GEN_35[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_sw = _GEN_35[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_sx = _GEN_35[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_sr = _GEN_35[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_pw = _GEN_35[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_px = _GEN_35[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_pr = _GEN_35[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_ppp = _GEN_35[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_pal = _GEN_35[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_paa = _GEN_35[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_eff = _GEN_35[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_c = _GEN_35[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_ppn = _GEN_39[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_u = _GEN_39[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_ae = _GEN_39[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_sw = _GEN_39[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_sx = _GEN_39[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_sr = _GEN_39[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_pw = _GEN_39[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_px = _GEN_39[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_pr = _GEN_39[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_ppp = _GEN_39[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_pal = _GEN_39[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_paa = _GEN_39[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_eff = _GEN_39[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_c = _GEN_39[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_ppn = _GEN_43[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_u = _GEN_43[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_ae = _GEN_43[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_sw = _GEN_43[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_sx = _GEN_43[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_sr = _GEN_43[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_pw = _GEN_43[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_px = _GEN_43[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_pr = _GEN_43[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_ppp = _GEN_43[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_pal = _GEN_43[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_paa = _GEN_43[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_eff = _GEN_43[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_c = _GEN_43[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_ppn = _GEN_47[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_u = _GEN_47[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_ae = _GEN_47[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_sw = _GEN_47[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_sx = _GEN_47[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_sr = _GEN_47[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_pw = _GEN_47[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_px = _GEN_47[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_pr = _GEN_47[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_ppp = _GEN_47[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_pal = _GEN_47[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_paa = _GEN_47[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_eff = _GEN_47[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_c = _GEN_47[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_ppn = _GEN_51[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_u = _GEN_51[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_ae = _GEN_51[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_sw = _GEN_51[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_sx = _GEN_51[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_sr = _GEN_51[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_pw = _GEN_51[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_px = _GEN_51[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_pr = _GEN_51[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_ppp = _GEN_51[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_pal = _GEN_51[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_paa = _GEN_51[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_eff = _GEN_51[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_c = _GEN_51[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_ppn = _GEN_55[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_u = _GEN_55[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_ae = _GEN_55[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_sw = _GEN_55[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_sx = _GEN_55[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_sr = _GEN_55[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_pw = _GEN_55[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_px = _GEN_55[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_pr = _GEN_55[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_ppp = _GEN_55[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_pal = _GEN_55[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_paa = _GEN_55[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_eff = _GEN_55[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_c = _GEN_55[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_ppn = _GEN_59[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_u = _GEN_59[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_ae = _GEN_59[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_sw = _GEN_59[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_sx = _GEN_59[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_sr = _GEN_59[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_pw = _GEN_59[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_px = _GEN_59[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_pr = _GEN_59[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_ppp = _GEN_59[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_pal = _GEN_59[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_paa = _GEN_59[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_eff = _GEN_59[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_c = _GEN_59[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_ppn = _GEN_63[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_u = _GEN_63[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_ae = _GEN_63[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_sw = _GEN_63[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_sx = _GEN_63[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_sr = _GEN_63[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_pw = _GEN_63[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_px = _GEN_63[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_pr = _GEN_63[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_ppp = _GEN_63[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_pal = _GEN_63[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_paa = _GEN_63[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_eff = _GEN_63[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_c = _GEN_63[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_u = superpage_entries_0_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_ae = superpage_entries_0_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_sw = superpage_entries_0_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_sx = superpage_entries_0_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_sr = superpage_entries_0_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_pw = superpage_entries_0_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_px = superpage_entries_0_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_pr = superpage_entries_0_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_ppp = superpage_entries_0_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_u = superpage_entries_1_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_ae = superpage_entries_1_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_sw = superpage_entries_1_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_sx = superpage_entries_1_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_sr = superpage_entries_1_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_pw = superpage_entries_1_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_px = superpage_entries_1_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_pr = superpage_entries_1_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_ppp = superpage_entries_1_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_u = superpage_entries_2_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_ae = superpage_entries_2_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_sw = superpage_entries_2_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_sx = superpage_entries_2_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_sr = superpage_entries_2_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_pw = superpage_entries_2_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_px = superpage_entries_2_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_pr = superpage_entries_2_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_ppp = superpage_entries_2_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_u = superpage_entries_3_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_ae = superpage_entries_3_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_sw = superpage_entries_3_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_sx = superpage_entries_3_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_sr = superpage_entries_3_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_pw = superpage_entries_3_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_px = superpage_entries_3_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_pr = superpage_entries_3_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_ppp = superpage_entries_3_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_u = special_entry_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_ae = special_entry_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_sw = special_entry_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_sx = special_entry_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_sr = special_entry_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_pw = special_entry_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_px = special_entry_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_pr = special_entry_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_ppp = special_entry_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_pal = special_entry_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_paa = special_entry_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_eff = special_entry_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_c = special_entry_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_ppn = _GEN_35[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_u = _GEN_35[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_ae = _GEN_35[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_sw = _GEN_35[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_sx = _GEN_35[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_sr = _GEN_35[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_pw = _GEN_35[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_px = _GEN_35[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_pr = _GEN_35[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_ppp = _GEN_35[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_pal = _GEN_35[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_paa = _GEN_35[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_eff = _GEN_35[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_c = _GEN_35[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_ppn = _GEN_39[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_u = _GEN_39[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_ae = _GEN_39[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_sw = _GEN_39[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_sx = _GEN_39[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_sr = _GEN_39[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_pw = _GEN_39[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_px = _GEN_39[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_pr = _GEN_39[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_ppp = _GEN_39[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_pal = _GEN_39[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_paa = _GEN_39[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_eff = _GEN_39[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_c = _GEN_39[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_ppn = _GEN_43[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_u = _GEN_43[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_ae = _GEN_43[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_sw = _GEN_43[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_sx = _GEN_43[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_sr = _GEN_43[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_pw = _GEN_43[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_px = _GEN_43[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_pr = _GEN_43[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_ppp = _GEN_43[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_pal = _GEN_43[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_paa = _GEN_43[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_eff = _GEN_43[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_c = _GEN_43[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_ppn = _GEN_47[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_u = _GEN_47[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_ae = _GEN_47[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_sw = _GEN_47[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_sx = _GEN_47[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_sr = _GEN_47[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_pw = _GEN_47[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_px = _GEN_47[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_pr = _GEN_47[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_ppp = _GEN_47[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_pal = _GEN_47[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_paa = _GEN_47[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_eff = _GEN_47[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_c = _GEN_47[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_ppn = _GEN_51[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_u = _GEN_51[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_ae = _GEN_51[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_sw = _GEN_51[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_sx = _GEN_51[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_sr = _GEN_51[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_pw = _GEN_51[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_px = _GEN_51[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_pr = _GEN_51[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_ppp = _GEN_51[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_pal = _GEN_51[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_paa = _GEN_51[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_eff = _GEN_51[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_c = _GEN_51[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_ppn = _GEN_55[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_u = _GEN_55[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_ae = _GEN_55[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_sw = _GEN_55[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_sx = _GEN_55[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_sr = _GEN_55[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_pw = _GEN_55[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_px = _GEN_55[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_pr = _GEN_55[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_ppp = _GEN_55[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_pal = _GEN_55[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_paa = _GEN_55[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_eff = _GEN_55[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_c = _GEN_55[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_ppn = _GEN_59[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_u = _GEN_59[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_ae = _GEN_59[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_sw = _GEN_59[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_sx = _GEN_59[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_sr = _GEN_59[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_pw = _GEN_59[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_px = _GEN_59[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_pr = _GEN_59[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_ppp = _GEN_59[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_pal = _GEN_59[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_paa = _GEN_59[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_eff = _GEN_59[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_c = _GEN_59[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_ppn = _GEN_63[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_u = _GEN_63[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_ae = _GEN_63[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_sw = _GEN_63[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_sx = _GEN_63[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_sr = _GEN_63[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_pw = _GEN_63[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_px = _GEN_63[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_pr = _GEN_63[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_ppp = _GEN_63[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_pal = _GEN_63[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_paa = _GEN_63[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_eff = _GEN_63[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_c = _GEN_63[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_u = superpage_entries_0_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_ae = superpage_entries_0_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_sw = superpage_entries_0_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_sx = superpage_entries_0_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_sr = superpage_entries_0_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_pw = superpage_entries_0_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_px = superpage_entries_0_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_pr = superpage_entries_0_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_ppp = superpage_entries_0_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_u = superpage_entries_1_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_ae = superpage_entries_1_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_sw = superpage_entries_1_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_sx = superpage_entries_1_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_sr = superpage_entries_1_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_pw = superpage_entries_1_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_px = superpage_entries_1_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_pr = superpage_entries_1_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_ppp = superpage_entries_1_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_u = superpage_entries_2_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_ae = superpage_entries_2_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_sw = superpage_entries_2_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_sx = superpage_entries_2_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_sr = superpage_entries_2_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_pw = superpage_entries_2_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_px = superpage_entries_2_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_pr = superpage_entries_2_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_ppp = superpage_entries_2_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_u = superpage_entries_3_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_ae = superpage_entries_3_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_sw = superpage_entries_3_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_sx = superpage_entries_3_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_sr = superpage_entries_3_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_pw = superpage_entries_3_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_px = superpage_entries_3_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_pr = superpage_entries_3_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_ppp = superpage_entries_3_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_u = special_entry_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_ae = special_entry_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_sw = special_entry_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_sx = special_entry_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_sr = special_entry_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_pw = special_entry_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_px = special_entry_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_pr = special_entry_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_ppp = special_entry_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_pal = special_entry_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_paa = special_entry_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_eff = special_entry_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_c = special_entry_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_ppn = _GEN_35[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_u = _GEN_35[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_ae = _GEN_35[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_sw = _GEN_35[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_sx = _GEN_35[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_sr = _GEN_35[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_pw = _GEN_35[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_px = _GEN_35[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_pr = _GEN_35[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_ppp = _GEN_35[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_pal = _GEN_35[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_paa = _GEN_35[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_eff = _GEN_35[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_c = _GEN_35[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_ppn = _GEN_39[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_u = _GEN_39[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_ae = _GEN_39[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_sw = _GEN_39[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_sx = _GEN_39[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_sr = _GEN_39[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_pw = _GEN_39[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_px = _GEN_39[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_pr = _GEN_39[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_ppp = _GEN_39[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_pal = _GEN_39[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_paa = _GEN_39[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_eff = _GEN_39[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_c = _GEN_39[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_ppn = _GEN_43[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_u = _GEN_43[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_ae = _GEN_43[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_sw = _GEN_43[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_sx = _GEN_43[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_sr = _GEN_43[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_pw = _GEN_43[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_px = _GEN_43[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_pr = _GEN_43[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_ppp = _GEN_43[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_pal = _GEN_43[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_paa = _GEN_43[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_eff = _GEN_43[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_c = _GEN_43[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_ppn = _GEN_47[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_u = _GEN_47[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_ae = _GEN_47[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_sw = _GEN_47[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_sx = _GEN_47[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_sr = _GEN_47[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_pw = _GEN_47[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_px = _GEN_47[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_pr = _GEN_47[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_ppp = _GEN_47[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_pal = _GEN_47[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_paa = _GEN_47[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_eff = _GEN_47[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_c = _GEN_47[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_ppn = _GEN_51[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_u = _GEN_51[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_ae = _GEN_51[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_sw = _GEN_51[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_sx = _GEN_51[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_sr = _GEN_51[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_pw = _GEN_51[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_px = _GEN_51[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_pr = _GEN_51[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_ppp = _GEN_51[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_pal = _GEN_51[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_paa = _GEN_51[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_eff = _GEN_51[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_c = _GEN_51[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_ppn = _GEN_55[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_u = _GEN_55[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_ae = _GEN_55[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_sw = _GEN_55[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_sx = _GEN_55[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_sr = _GEN_55[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_pw = _GEN_55[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_px = _GEN_55[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_pr = _GEN_55[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_ppp = _GEN_55[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_pal = _GEN_55[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_paa = _GEN_55[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_eff = _GEN_55[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_c = _GEN_55[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_ppn = _GEN_59[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_u = _GEN_59[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_ae = _GEN_59[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_sw = _GEN_59[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_sx = _GEN_59[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_sr = _GEN_59[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_pw = _GEN_59[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_px = _GEN_59[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_pr = _GEN_59[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_ppp = _GEN_59[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_pal = _GEN_59[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_paa = _GEN_59[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_eff = _GEN_59[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_c = _GEN_59[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_ppn = _GEN_63[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_u = _GEN_63[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_ae = _GEN_63[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_sw = _GEN_63[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_sx = _GEN_63[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_sr = _GEN_63[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_pw = _GEN_63[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_px = _GEN_63[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_pr = _GEN_63[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_ppp = _GEN_63[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_pal = _GEN_63[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_paa = _GEN_63[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_eff = _GEN_63[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_c = _GEN_63[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_u = superpage_entries_0_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_ae = superpage_entries_0_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_sw = superpage_entries_0_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_sx = superpage_entries_0_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_sr = superpage_entries_0_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_pw = superpage_entries_0_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_px = superpage_entries_0_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_pr = superpage_entries_0_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_ppp = superpage_entries_0_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_u = superpage_entries_1_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_ae = superpage_entries_1_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_sw = superpage_entries_1_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_sx = superpage_entries_1_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_sr = superpage_entries_1_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_pw = superpage_entries_1_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_px = superpage_entries_1_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_pr = superpage_entries_1_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_ppp = superpage_entries_1_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_u = superpage_entries_2_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_ae = superpage_entries_2_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_sw = superpage_entries_2_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_sx = superpage_entries_2_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_sr = superpage_entries_2_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_pw = superpage_entries_2_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_px = superpage_entries_2_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_pr = superpage_entries_2_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_ppp = superpage_entries_2_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_u = superpage_entries_3_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_ae = superpage_entries_3_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_sw = superpage_entries_3_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_sx = superpage_entries_3_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_sr = superpage_entries_3_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_pw = superpage_entries_3_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_px = superpage_entries_3_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_pr = superpage_entries_3_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_ppp = superpage_entries_3_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 244:18]
  assign TLB_cov_read_addr = TLB_state;
  assign TLB_cov_read_data = TLB_cov[TLB_cov_read_addr]; // @[Coverage map for TLB]
  assign TLB_cov_write_data = 1'h1;
  assign TLB_cov_write_addr = TLB_state;
  assign TLB_cov_write_mask = 1'h1;
  assign TLB_cov_write_en = 1'h1;
  assign mux_cond_0 = sectored_entries_7_data_2[0];
  assign mux_cond_1 = ~sectored_entries_1_data_1[13];
  assign mux_cond_2 = ~sectored_entries_4_data_3[13];
  assign mux_cond_3 = ~sectored_entries_3_data_3[13];
  assign mux_cond_4 = sectored_entries_4_data_0[0];
  assign mux_cond_5 = sectored_entries_0_data_1[0];
  assign mux_cond_6 = sectored_entries_0_data_0[0];
  assign mux_cond_7 = sectored_entries_4_data_3[0];
  assign mux_cond_8 = sectored_entries_1_data_3[0];
  assign mux_cond_9 = sectored_entries_2_data_1[0];
  assign mux_cond_10 = ~sectored_entries_6_data_1[13];
  assign mux_cond_11 = ~sectored_entries_1_data_0[13];
  assign mux_cond_12 = sectored_entries_6_data_2[0];
  assign mux_cond_13 = ~sectored_entries_4_data_1[13];
  assign mux_cond_14 = sectored_entries_6_data_0[0];
  assign mux_cond_15 = sectored_entries_7_data_0[0];
  assign mux_cond_16 = sectored_entries_2_data_2[0];
  assign mux_cond_17 = sectored_entries_7_data_3[0];
  assign mux_cond_18 = ~sectored_entries_2_data_1[13];
  assign mux_cond_19 = sectored_entries_4_data_2[0];
  assign mux_cond_20 = ~sectored_entries_1_data_2[13];
  assign mux_cond_21 = ~superpage_entries_1_data_0[13];
  assign mux_cond_22 = ~sectored_entries_2_data_2[13];
  assign mux_cond_23 = ~sectored_entries_7_data_2[13];
  assign mux_cond_24 = ~sectored_entries_6_data_2[13];
  assign mux_cond_25 = ~sectored_entries_3_data_0[13];
  assign mux_cond_26 = sectored_entries_5_data_1[0];
  assign mux_cond_27 = sectored_entries_5_data_3[0];
  assign mux_cond_28 = ~sectored_entries_5_data_2[13];
  assign mux_cond_29 = sectored_entries_6_data_3[0];
  assign mux_cond_30 = ~sectored_entries_3_data_2[13];
  assign mux_cond_31 = ~sectored_entries_3_data_1[13];
  assign mux_cond_32 = sectored_entries_3_data_2[0];
  assign mux_cond_33 = ~sectored_entries_6_data_0[13];
  assign mux_cond_34 = sectored_entries_1_data_1[0];
  assign mux_cond_35 = ~sectored_entries_0_data_1[13];
  assign mux_cond_36 = sectored_entries_6_data_1[0];
  assign mux_cond_37 = sectored_entries_3_data_3[0];
  assign mux_cond_38 = ~sectored_entries_0_data_0[13];
  assign mux_cond_39 = sectored_entries_1_data_0[0];
  assign mux_cond_40 = ~sectored_entries_2_data_3[13];
  assign mux_cond_41 = sectored_entries_5_data_2[0];
  assign mux_cond_42 = sectored_entries_7_data_1[0];
  assign mux_cond_43 = ~sectored_entries_7_data_1[13];
  assign mux_cond_44 = sectored_entries_0_data_2[0];
  assign mux_cond_45 = sectored_entries_0_data_3[0];
  assign mux_cond_46 = ~sectored_entries_6_data_3[13];
  assign mux_cond_47 = sectored_entries_3_data_0[0];
  assign mux_cond_48 = ~sectored_entries_0_data_3[13];
  assign mux_cond_49 = sectored_entries_1_data_2[0];
  assign mux_cond_50 = sectored_entries_2_data_3[0];
  assign mux_cond_51 = sectored_entries_5_data_0[0];
  assign mux_cond_52 = ~sectored_entries_5_data_1[13];
  assign mux_cond_53 = ~sectored_entries_2_data_0[13];
  assign mux_cond_54 = ~sectored_entries_7_data_0[13];
  assign mux_cond_55 = ~sectored_entries_5_data_0[13];
  assign mux_cond_56 = ~sectored_entries_0_data_2[13];
  assign mux_cond_57 = ~superpage_entries_3_data_0[13];
  assign mux_cond_58 = ~special_entry_data_0[13];
  assign mux_cond_59 = sectored_entries_3_data_1[0];
  assign mux_cond_60 = sectored_entries_2_data_0[0];
  assign mux_cond_61 = ~sectored_entries_4_data_2[13];
  assign mux_cond_62 = ~sectored_entries_1_data_3[13];
  assign mux_cond_63 = ~superpage_entries_0_data_0[13];
  assign mux_cond_64 = sectored_entries_4_data_1[0];
  assign mux_cond_65 = ~sectored_entries_5_data_3[13];
  assign mux_cond_66 = ~superpage_entries_2_data_0[13];
  assign mux_cond_67 = ~sectored_entries_4_data_0[13];
  assign mux_cond_68 = ~sectored_entries_7_data_3[13];
  assign state_shl = {state, 5'h0};
  assign state_pad = {13'h0,state_shl};
  assign r_sectored_repl_addr_shl = {r_sectored_repl_addr, 12'h0};
  assign r_sectored_repl_addr_pad = {5'h0,r_sectored_repl_addr_shl};
  assign r_superpage_repl_addr_shl = {r_superpage_repl_addr, 2'h0};
  assign r_superpage_repl_addr_pad = {16'h0,r_superpage_repl_addr_shl};
  assign r_sectored_hit_addr_shl = {r_sectored_hit_addr, 8'h0};
  assign r_sectored_hit_addr_pad = {9'h0,r_sectored_hit_addr_shl};
  assign special_entry_valid_0_shl = {special_entry_valid_0, 15'h0};
  assign special_entry_valid_0_pad = {4'h0,special_entry_valid_0_shl};
  assign r_sectored_hit_shl = {r_sectored_hit, 12'h0};
  assign r_sectored_hit_pad = {7'h0,r_sectored_hit_shl};
  assign special_entry_level_shl = {special_entry_level, 3'h0};
  assign special_entry_level_pad = {15'h0,special_entry_level_shl};
  assign mux_cond_0_shl = {mux_cond_0, 8'h0};
  assign mux_cond_0_pad = {11'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 12'h0};
  assign mux_cond_1_pad = {7'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 5'h0};
  assign mux_cond_2_pad = {14'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 7'h0};
  assign mux_cond_3_pad = {12'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 7'h0};
  assign mux_cond_4_pad = {12'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 5'h0};
  assign mux_cond_5_pad = {14'h0,mux_cond_5_shl};
  assign mux_cond_6_shl = {mux_cond_6, 4'h0};
  assign mux_cond_6_pad = {15'h0,mux_cond_6_shl};
  assign mux_cond_7_shl = {mux_cond_7, 18'h0};
  assign mux_cond_7_pad = {1'h0,mux_cond_7_shl};
  assign mux_cond_8_shl = {mux_cond_8, 2'h0};
  assign mux_cond_8_pad = {17'h0,mux_cond_8_shl};
  assign mux_cond_9_shl = {mux_cond_9, 6'h0};
  assign mux_cond_9_pad = {13'h0,mux_cond_9_shl};
  assign mux_cond_10_shl = mux_cond_10;
  assign mux_cond_10_pad = {19'h0,mux_cond_10_shl};
  assign mux_cond_11_shl = {mux_cond_11, 14'h0};
  assign mux_cond_11_pad = {5'h0,mux_cond_11_shl};
  assign mux_cond_12_shl = {mux_cond_12, 15'h0};
  assign mux_cond_12_pad = {4'h0,mux_cond_12_shl};
  assign mux_cond_13_shl = mux_cond_13;
  assign mux_cond_13_pad = {19'h0,mux_cond_13_shl};
  assign mux_cond_14_shl = {mux_cond_14, 17'h0};
  assign mux_cond_14_pad = {2'h0,mux_cond_14_shl};
  assign mux_cond_15_shl = {mux_cond_15, 9'h0};
  assign mux_cond_15_pad = {10'h0,mux_cond_15_shl};
  assign mux_cond_16_shl = {mux_cond_16, 4'h0};
  assign mux_cond_16_pad = {15'h0,mux_cond_16_shl};
  assign mux_cond_17_shl = {mux_cond_17, 7'h0};
  assign mux_cond_17_pad = {12'h0,mux_cond_17_shl};
  assign mux_cond_18_shl = {mux_cond_18, 15'h0};
  assign mux_cond_18_pad = {4'h0,mux_cond_18_shl};
  assign mux_cond_19_shl = {mux_cond_19, 10'h0};
  assign mux_cond_19_pad = {9'h0,mux_cond_19_shl};
  assign mux_cond_20_shl = {mux_cond_20, 4'h0};
  assign mux_cond_20_pad = {15'h0,mux_cond_20_shl};
  assign mux_cond_21_shl = {mux_cond_21, 5'h0};
  assign mux_cond_21_pad = {14'h0,mux_cond_21_shl};
  assign mux_cond_22_shl = {mux_cond_22, 7'h0};
  assign mux_cond_22_pad = {12'h0,mux_cond_22_shl};
  assign mux_cond_23_shl = {mux_cond_23, 17'h0};
  assign mux_cond_23_pad = {2'h0,mux_cond_23_shl};
  assign mux_cond_24_shl = {mux_cond_24, 8'h0};
  assign mux_cond_24_pad = {11'h0,mux_cond_24_shl};
  assign mux_cond_25_shl = {mux_cond_25, 7'h0};
  assign mux_cond_25_pad = {12'h0,mux_cond_25_shl};
  assign mux_cond_26_shl = {mux_cond_26, 18'h0};
  assign mux_cond_26_pad = {1'h0,mux_cond_26_shl};
  assign mux_cond_27_shl = {mux_cond_27, 9'h0};
  assign mux_cond_27_pad = {10'h0,mux_cond_27_shl};
  assign mux_cond_28_shl = {mux_cond_28, 10'h0};
  assign mux_cond_28_pad = {9'h0,mux_cond_28_shl};
  assign mux_cond_29_shl = {mux_cond_29, 9'h0};
  assign mux_cond_29_pad = {10'h0,mux_cond_29_shl};
  assign mux_cond_30_shl = {mux_cond_30, 16'h0};
  assign mux_cond_30_pad = {3'h0,mux_cond_30_shl};
  assign mux_cond_31_shl = {mux_cond_31, 3'h0};
  assign mux_cond_31_pad = {16'h0,mux_cond_31_shl};
  assign mux_cond_32_shl = {mux_cond_32, 1'h0};
  assign mux_cond_32_pad = {18'h0,mux_cond_32_shl};
  assign mux_cond_33_shl = {mux_cond_33, 5'h0};
  assign mux_cond_33_pad = {14'h0,mux_cond_33_shl};
  assign mux_cond_34_shl = {mux_cond_34, 4'h0};
  assign mux_cond_34_pad = {15'h0,mux_cond_34_shl};
  assign mux_cond_35_shl = {mux_cond_35, 12'h0};
  assign mux_cond_35_pad = {7'h0,mux_cond_35_shl};
  assign mux_cond_36_shl = {mux_cond_36, 9'h0};
  assign mux_cond_36_pad = {10'h0,mux_cond_36_shl};
  assign mux_cond_37_shl = {mux_cond_37, 4'h0};
  assign mux_cond_37_pad = {15'h0,mux_cond_37_shl};
  assign mux_cond_38_shl = {mux_cond_38, 10'h0};
  assign mux_cond_38_pad = {9'h0,mux_cond_38_shl};
  assign mux_cond_39_shl = {mux_cond_39, 8'h0};
  assign mux_cond_39_pad = {11'h0,mux_cond_39_shl};
  assign mux_cond_40_shl = {mux_cond_40, 18'h0};
  assign mux_cond_40_pad = {1'h0,mux_cond_40_shl};
  assign mux_cond_41_shl = {mux_cond_41, 17'h0};
  assign mux_cond_41_pad = {2'h0,mux_cond_41_shl};
  assign mux_cond_42_shl = {mux_cond_42, 18'h0};
  assign mux_cond_42_pad = {1'h0,mux_cond_42_shl};
  assign mux_cond_43_shl = {mux_cond_43, 18'h0};
  assign mux_cond_43_pad = {1'h0,mux_cond_43_shl};
  assign mux_cond_44_shl = mux_cond_44;
  assign mux_cond_44_pad = {19'h0,mux_cond_44_shl};
  assign mux_cond_45_shl = {mux_cond_45, 11'h0};
  assign mux_cond_45_pad = {8'h0,mux_cond_45_shl};
  assign mux_cond_46_shl = {mux_cond_46, 15'h0};
  assign mux_cond_46_pad = {4'h0,mux_cond_46_shl};
  assign mux_cond_47_shl = {mux_cond_47, 6'h0};
  assign mux_cond_47_pad = {13'h0,mux_cond_47_shl};
  assign mux_cond_48_shl = mux_cond_48;
  assign mux_cond_48_pad = {19'h0,mux_cond_48_shl};
  assign mux_cond_49_shl = {mux_cond_49, 18'h0};
  assign mux_cond_49_pad = {1'h0,mux_cond_49_shl};
  assign mux_cond_50_shl = {mux_cond_50, 19'h0};
  assign mux_cond_50_pad = mux_cond_50_shl;
  assign mux_cond_51_shl = {mux_cond_51, 7'h0};
  assign mux_cond_51_pad = {12'h0,mux_cond_51_shl};
  assign mux_cond_52_shl = {mux_cond_52, 18'h0};
  assign mux_cond_52_pad = {1'h0,mux_cond_52_shl};
  assign mux_cond_53_shl = {mux_cond_53, 17'h0};
  assign mux_cond_53_pad = {2'h0,mux_cond_53_shl};
  assign mux_cond_54_shl = {mux_cond_54, 17'h0};
  assign mux_cond_54_pad = {2'h0,mux_cond_54_shl};
  assign mux_cond_55_shl = {mux_cond_55, 15'h0};
  assign mux_cond_55_pad = {4'h0,mux_cond_55_shl};
  assign mux_cond_56_shl = {mux_cond_56, 4'h0};
  assign mux_cond_56_pad = {15'h0,mux_cond_56_shl};
  assign mux_cond_57_shl = {mux_cond_57, 3'h0};
  assign mux_cond_57_pad = {16'h0,mux_cond_57_shl};
  assign mux_cond_58_shl = {mux_cond_58, 6'h0};
  assign mux_cond_58_pad = {13'h0,mux_cond_58_shl};
  assign mux_cond_59_shl = {mux_cond_59, 10'h0};
  assign mux_cond_59_pad = {9'h0,mux_cond_59_shl};
  assign mux_cond_60_shl = {mux_cond_60, 15'h0};
  assign mux_cond_60_pad = {4'h0,mux_cond_60_shl};
  assign mux_cond_61_shl = {mux_cond_61, 19'h0};
  assign mux_cond_61_pad = mux_cond_61_shl;
  assign mux_cond_62_shl = {mux_cond_62, 14'h0};
  assign mux_cond_62_pad = {5'h0,mux_cond_62_shl};
  assign mux_cond_63_shl = {mux_cond_63, 11'h0};
  assign mux_cond_63_pad = {8'h0,mux_cond_63_shl};
  assign mux_cond_64_shl = {mux_cond_64, 2'h0};
  assign mux_cond_64_pad = {17'h0,mux_cond_64_shl};
  assign mux_cond_65_shl = {mux_cond_65, 7'h0};
  assign mux_cond_65_pad = {12'h0,mux_cond_65_shl};
  assign mux_cond_66_shl = {mux_cond_66, 3'h0};
  assign mux_cond_66_pad = {16'h0,mux_cond_66_shl};
  assign mux_cond_67_shl = {mux_cond_67, 1'h0};
  assign mux_cond_67_pad = {18'h0,mux_cond_67_shl};
  assign mux_cond_68_shl = {mux_cond_68, 7'h0};
  assign mux_cond_68_pad = {12'h0,mux_cond_68_shl};
  assign superpage_entries_2_level_shl = {superpage_entries_2_level, 18'h0};
  assign superpage_entries_2_level_pad = superpage_entries_2_level_shl;
  assign sectored_entries_7_valid_3_shl = {sectored_entries_7_valid_3, 2'h0};
  assign sectored_entries_7_valid_3_pad = {17'h0,sectored_entries_7_valid_3_shl};
  assign superpage_entries_1_level_shl = {superpage_entries_1_level, 18'h0};
  assign superpage_entries_1_level_pad = superpage_entries_1_level_shl;
  assign superpage_entries_1_valid_0_shl = {superpage_entries_1_valid_0, 18'h0};
  assign superpage_entries_1_valid_0_pad = {1'h0,superpage_entries_1_valid_0_shl};
  assign sectored_entries_3_valid_0_shl = {sectored_entries_3_valid_0, 10'h0};
  assign sectored_entries_3_valid_0_pad = {9'h0,sectored_entries_3_valid_0_shl};
  assign sectored_entries_1_valid_3_shl = {sectored_entries_1_valid_3, 2'h0};
  assign sectored_entries_1_valid_3_pad = {17'h0,sectored_entries_1_valid_3_shl};
  assign sectored_entries_6_valid_3_shl = {sectored_entries_6_valid_3, 2'h0};
  assign sectored_entries_6_valid_3_pad = {17'h0,sectored_entries_6_valid_3_shl};
  assign sectored_entries_1_valid_0_shl = {sectored_entries_1_valid_0, 10'h0};
  assign sectored_entries_1_valid_0_pad = {9'h0,sectored_entries_1_valid_0_shl};
  assign sectored_entries_2_valid_0_shl = {sectored_entries_2_valid_0, 10'h0};
  assign sectored_entries_2_valid_0_pad = {9'h0,sectored_entries_2_valid_0_shl};
  assign sectored_entries_3_valid_1_shl = {sectored_entries_3_valid_1, 5'h0};
  assign sectored_entries_3_valid_1_pad = {14'h0,sectored_entries_3_valid_1_shl};
  assign sectored_entries_5_valid_3_shl = {sectored_entries_5_valid_3, 2'h0};
  assign sectored_entries_5_valid_3_pad = {17'h0,sectored_entries_5_valid_3_shl};
  assign superpage_entries_3_valid_0_shl = {superpage_entries_3_valid_0, 18'h0};
  assign superpage_entries_3_valid_0_pad = {1'h0,superpage_entries_3_valid_0_shl};
  assign sectored_entries_5_valid_1_shl = {sectored_entries_5_valid_1, 5'h0};
  assign sectored_entries_5_valid_1_pad = {14'h0,sectored_entries_5_valid_1_shl};
  assign sectored_entries_0_valid_3_shl = {sectored_entries_0_valid_3, 2'h0};
  assign sectored_entries_0_valid_3_pad = {17'h0,sectored_entries_0_valid_3_shl};
  assign sectored_entries_6_valid_0_shl = {sectored_entries_6_valid_0, 10'h0};
  assign sectored_entries_6_valid_0_pad = {9'h0,sectored_entries_6_valid_0_shl};
  assign sectored_entries_0_valid_0_shl = {sectored_entries_0_valid_0, 10'h0};
  assign sectored_entries_0_valid_0_pad = {9'h0,sectored_entries_0_valid_0_shl};
  assign sectored_entries_4_valid_2_shl = {sectored_entries_4_valid_2, 5'h0};
  assign sectored_entries_4_valid_2_pad = {14'h0,sectored_entries_4_valid_2_shl};
  assign superpage_entries_2_valid_0_shl = {superpage_entries_2_valid_0, 18'h0};
  assign superpage_entries_2_valid_0_pad = {1'h0,superpage_entries_2_valid_0_shl};
  assign sectored_entries_2_valid_1_shl = {sectored_entries_2_valid_1, 5'h0};
  assign sectored_entries_2_valid_1_pad = {14'h0,sectored_entries_2_valid_1_shl};
  assign superpage_entries_0_level_shl = {superpage_entries_0_level, 18'h0};
  assign superpage_entries_0_level_pad = superpage_entries_0_level_shl;
  assign sectored_entries_1_valid_1_shl = {sectored_entries_1_valid_1, 5'h0};
  assign sectored_entries_1_valid_1_pad = {14'h0,sectored_entries_1_valid_1_shl};
  assign sectored_entries_4_valid_3_shl = {sectored_entries_4_valid_3, 2'h0};
  assign sectored_entries_4_valid_3_pad = {17'h0,sectored_entries_4_valid_3_shl};
  assign sectored_entries_0_valid_1_shl = {sectored_entries_0_valid_1, 5'h0};
  assign sectored_entries_0_valid_1_pad = {14'h0,sectored_entries_0_valid_1_shl};
  assign sectored_entries_4_valid_0_shl = {sectored_entries_4_valid_0, 10'h0};
  assign sectored_entries_4_valid_0_pad = {9'h0,sectored_entries_4_valid_0_shl};
  assign sectored_entries_0_valid_2_shl = {sectored_entries_0_valid_2, 5'h0};
  assign sectored_entries_0_valid_2_pad = {14'h0,sectored_entries_0_valid_2_shl};
  assign sectored_entries_1_valid_2_shl = {sectored_entries_1_valid_2, 5'h0};
  assign sectored_entries_1_valid_2_pad = {14'h0,sectored_entries_1_valid_2_shl};
  assign sectored_entries_2_valid_2_shl = {sectored_entries_2_valid_2, 5'h0};
  assign sectored_entries_2_valid_2_pad = {14'h0,sectored_entries_2_valid_2_shl};
  assign sectored_entries_7_valid_0_shl = {sectored_entries_7_valid_0, 10'h0};
  assign sectored_entries_7_valid_0_pad = {9'h0,sectored_entries_7_valid_0_shl};
  assign sectored_entries_5_valid_2_shl = {sectored_entries_5_valid_2, 5'h0};
  assign sectored_entries_5_valid_2_pad = {14'h0,sectored_entries_5_valid_2_shl};
  assign sectored_entries_7_valid_2_shl = {sectored_entries_7_valid_2, 5'h0};
  assign sectored_entries_7_valid_2_pad = {14'h0,sectored_entries_7_valid_2_shl};
  assign sectored_entries_4_valid_1_shl = {sectored_entries_4_valid_1, 5'h0};
  assign sectored_entries_4_valid_1_pad = {14'h0,sectored_entries_4_valid_1_shl};
  assign sectored_entries_5_valid_0_shl = {sectored_entries_5_valid_0, 10'h0};
  assign sectored_entries_5_valid_0_pad = {9'h0,sectored_entries_5_valid_0_shl};
  assign sectored_entries_7_valid_1_shl = {sectored_entries_7_valid_1, 5'h0};
  assign sectored_entries_7_valid_1_pad = {14'h0,sectored_entries_7_valid_1_shl};
  assign superpage_entries_3_level_shl = {superpage_entries_3_level, 18'h0};
  assign superpage_entries_3_level_pad = superpage_entries_3_level_shl;
  assign sectored_entries_3_valid_3_shl = {sectored_entries_3_valid_3, 2'h0};
  assign sectored_entries_3_valid_3_pad = {17'h0,sectored_entries_3_valid_3_shl};
  assign sectored_entries_2_valid_3_shl = {sectored_entries_2_valid_3, 2'h0};
  assign sectored_entries_2_valid_3_pad = {17'h0,sectored_entries_2_valid_3_shl};
  assign superpage_entries_0_valid_0_shl = {superpage_entries_0_valid_0, 18'h0};
  assign superpage_entries_0_valid_0_pad = {1'h0,superpage_entries_0_valid_0_shl};
  assign sectored_entries_6_valid_1_shl = {sectored_entries_6_valid_1, 5'h0};
  assign sectored_entries_6_valid_1_pad = {14'h0,sectored_entries_6_valid_1_shl};
  assign sectored_entries_3_valid_2_shl = {sectored_entries_3_valid_2, 5'h0};
  assign sectored_entries_3_valid_2_pad = {14'h0,sectored_entries_3_valid_2_shl};
  assign sectored_entries_6_valid_2_shl = {sectored_entries_6_valid_2, 5'h0};
  assign sectored_entries_6_valid_2_pad = {14'h0,sectored_entries_6_valid_2_shl};
  assign TLB_xor64 = r_sectored_repl_addr_pad ^ r_superpage_repl_addr_pad;
  assign TLB_xor31 = state_pad ^ TLB_xor64;
  assign TLB_xor65 = r_sectored_hit_addr_pad ^ special_entry_valid_0_pad;
  assign TLB_xor66 = r_sectored_hit_pad ^ special_entry_level_pad;
  assign TLB_xor32 = TLB_xor65 ^ TLB_xor66;
  assign TLB_xor15 = TLB_xor31 ^ TLB_xor32;
  assign TLB_xor68 = mux_cond_1_pad ^ mux_cond_2_pad;
  assign TLB_xor33 = mux_cond_0_pad ^ TLB_xor68;
  assign TLB_xor69 = mux_cond_3_pad ^ mux_cond_4_pad;
  assign TLB_xor70 = mux_cond_5_pad ^ mux_cond_6_pad;
  assign TLB_xor34 = TLB_xor69 ^ TLB_xor70;
  assign TLB_xor16 = TLB_xor33 ^ TLB_xor34;
  assign TLB_xor7 = TLB_xor15 ^ TLB_xor16;
  assign TLB_xor72 = mux_cond_8_pad ^ mux_cond_9_pad;
  assign TLB_xor35 = mux_cond_7_pad ^ TLB_xor72;
  assign TLB_xor73 = mux_cond_10_pad ^ mux_cond_11_pad;
  assign TLB_xor74 = mux_cond_12_pad ^ mux_cond_13_pad;
  assign TLB_xor36 = TLB_xor73 ^ TLB_xor74;
  assign TLB_xor17 = TLB_xor35 ^ TLB_xor36;
  assign TLB_xor75 = mux_cond_14_pad ^ mux_cond_15_pad;
  assign TLB_xor76 = mux_cond_16_pad ^ mux_cond_17_pad;
  assign TLB_xor37 = TLB_xor75 ^ TLB_xor76;
  assign TLB_xor77 = mux_cond_18_pad ^ mux_cond_19_pad;
  assign TLB_xor78 = mux_cond_20_pad ^ mux_cond_21_pad;
  assign TLB_xor38 = TLB_xor77 ^ TLB_xor78;
  assign TLB_xor18 = TLB_xor37 ^ TLB_xor38;
  assign TLB_xor8 = TLB_xor17 ^ TLB_xor18;
  assign TLB_xor3 = TLB_xor7 ^ TLB_xor8;
  assign TLB_xor80 = mux_cond_23_pad ^ mux_cond_24_pad;
  assign TLB_xor39 = mux_cond_22_pad ^ TLB_xor80;
  assign TLB_xor81 = mux_cond_25_pad ^ mux_cond_26_pad;
  assign TLB_xor82 = mux_cond_27_pad ^ mux_cond_28_pad;
  assign TLB_xor40 = TLB_xor81 ^ TLB_xor82;
  assign TLB_xor19 = TLB_xor39 ^ TLB_xor40;
  assign TLB_xor84 = mux_cond_30_pad ^ mux_cond_31_pad;
  assign TLB_xor41 = mux_cond_29_pad ^ TLB_xor84;
  assign TLB_xor85 = mux_cond_32_pad ^ mux_cond_33_pad;
  assign TLB_xor86 = mux_cond_34_pad ^ mux_cond_35_pad;
  assign TLB_xor42 = TLB_xor85 ^ TLB_xor86;
  assign TLB_xor20 = TLB_xor41 ^ TLB_xor42;
  assign TLB_xor9 = TLB_xor19 ^ TLB_xor20;
  assign TLB_xor88 = mux_cond_37_pad ^ mux_cond_38_pad;
  assign TLB_xor43 = mux_cond_36_pad ^ TLB_xor88;
  assign TLB_xor89 = mux_cond_39_pad ^ mux_cond_40_pad;
  assign TLB_xor90 = mux_cond_41_pad ^ mux_cond_42_pad;
  assign TLB_xor44 = TLB_xor89 ^ TLB_xor90;
  assign TLB_xor21 = TLB_xor43 ^ TLB_xor44;
  assign TLB_xor91 = mux_cond_43_pad ^ mux_cond_44_pad;
  assign TLB_xor92 = mux_cond_45_pad ^ mux_cond_46_pad;
  assign TLB_xor45 = TLB_xor91 ^ TLB_xor92;
  assign TLB_xor93 = mux_cond_47_pad ^ mux_cond_48_pad;
  assign TLB_xor94 = mux_cond_49_pad ^ mux_cond_50_pad;
  assign TLB_xor46 = TLB_xor93 ^ TLB_xor94;
  assign TLB_xor22 = TLB_xor45 ^ TLB_xor46;
  assign TLB_xor10 = TLB_xor21 ^ TLB_xor22;
  assign TLB_xor4 = TLB_xor9 ^ TLB_xor10;
  assign TLB_xor1 = TLB_xor3 ^ TLB_xor4;
  assign TLB_xor96 = mux_cond_52_pad ^ mux_cond_53_pad;
  assign TLB_xor47 = mux_cond_51_pad ^ TLB_xor96;
  assign TLB_xor97 = mux_cond_54_pad ^ mux_cond_55_pad;
  assign TLB_xor98 = mux_cond_56_pad ^ mux_cond_57_pad;
  assign TLB_xor48 = TLB_xor97 ^ TLB_xor98;
  assign TLB_xor23 = TLB_xor47 ^ TLB_xor48;
  assign TLB_xor100 = mux_cond_59_pad ^ mux_cond_60_pad;
  assign TLB_xor49 = mux_cond_58_pad ^ TLB_xor100;
  assign TLB_xor101 = mux_cond_61_pad ^ mux_cond_62_pad;
  assign TLB_xor102 = mux_cond_63_pad ^ mux_cond_64_pad;
  assign TLB_xor50 = TLB_xor101 ^ TLB_xor102;
  assign TLB_xor24 = TLB_xor49 ^ TLB_xor50;
  assign TLB_xor11 = TLB_xor23 ^ TLB_xor24;
  assign TLB_xor104 = mux_cond_66_pad ^ mux_cond_67_pad;
  assign TLB_xor51 = mux_cond_65_pad ^ TLB_xor104;
  assign TLB_xor105 = mux_cond_68_pad ^ superpage_entries_2_level_pad;
  assign TLB_xor106 = sectored_entries_7_valid_3_pad ^ superpage_entries_1_level_pad;
  assign TLB_xor52 = TLB_xor105 ^ TLB_xor106;
  assign TLB_xor25 = TLB_xor51 ^ TLB_xor52;
  assign TLB_xor107 = superpage_entries_1_valid_0_pad ^ sectored_entries_3_valid_0_pad;
  assign TLB_xor108 = sectored_entries_1_valid_3_pad ^ sectored_entries_6_valid_3_pad;
  assign TLB_xor53 = TLB_xor107 ^ TLB_xor108;
  assign TLB_xor109 = sectored_entries_1_valid_0_pad ^ sectored_entries_2_valid_0_pad;
  assign TLB_xor110 = sectored_entries_3_valid_1_pad ^ sectored_entries_5_valid_3_pad;
  assign TLB_xor54 = TLB_xor109 ^ TLB_xor110;
  assign TLB_xor26 = TLB_xor53 ^ TLB_xor54;
  assign TLB_xor12 = TLB_xor25 ^ TLB_xor26;
  assign TLB_xor5 = TLB_xor11 ^ TLB_xor12;
  assign TLB_xor112 = sectored_entries_5_valid_1_pad ^ sectored_entries_0_valid_3_pad;
  assign TLB_xor55 = superpage_entries_3_valid_0_pad ^ TLB_xor112;
  assign TLB_xor113 = sectored_entries_6_valid_0_pad ^ sectored_entries_0_valid_0_pad;
  assign TLB_xor114 = sectored_entries_4_valid_2_pad ^ superpage_entries_2_valid_0_pad;
  assign TLB_xor56 = TLB_xor113 ^ TLB_xor114;
  assign TLB_xor27 = TLB_xor55 ^ TLB_xor56;
  assign TLB_xor116 = superpage_entries_0_level_pad ^ sectored_entries_1_valid_1_pad;
  assign TLB_xor57 = sectored_entries_2_valid_1_pad ^ TLB_xor116;
  assign TLB_xor117 = sectored_entries_4_valid_3_pad ^ sectored_entries_0_valid_1_pad;
  assign TLB_xor118 = sectored_entries_4_valid_0_pad ^ sectored_entries_0_valid_2_pad;
  assign TLB_xor58 = TLB_xor117 ^ TLB_xor118;
  assign TLB_xor28 = TLB_xor57 ^ TLB_xor58;
  assign TLB_xor13 = TLB_xor27 ^ TLB_xor28;
  assign TLB_xor120 = sectored_entries_2_valid_2_pad ^ sectored_entries_7_valid_0_pad;
  assign TLB_xor59 = sectored_entries_1_valid_2_pad ^ TLB_xor120;
  assign TLB_xor121 = sectored_entries_5_valid_2_pad ^ sectored_entries_7_valid_2_pad;
  assign TLB_xor122 = sectored_entries_4_valid_1_pad ^ sectored_entries_5_valid_0_pad;
  assign TLB_xor60 = TLB_xor121 ^ TLB_xor122;
  assign TLB_xor29 = TLB_xor59 ^ TLB_xor60;
  assign TLB_xor123 = sectored_entries_7_valid_1_pad ^ superpage_entries_3_level_pad;
  assign TLB_xor124 = sectored_entries_3_valid_3_pad ^ sectored_entries_2_valid_3_pad;
  assign TLB_xor61 = TLB_xor123 ^ TLB_xor124;
  assign TLB_xor125 = superpage_entries_0_valid_0_pad ^ sectored_entries_6_valid_1_pad;
  assign TLB_xor126 = sectored_entries_3_valid_2_pad ^ sectored_entries_6_valid_2_pad;
  assign TLB_xor62 = TLB_xor125 ^ TLB_xor126;
  assign TLB_xor30 = TLB_xor61 ^ TLB_xor62;
  assign TLB_xor14 = TLB_xor29 ^ TLB_xor30;
  assign TLB_xor6 = TLB_xor13 ^ TLB_xor14;
  assign TLB_xor2 = TLB_xor5 ^ TLB_xor6;
  assign TLB_xor0 = TLB_xor1 ^ TLB_xor2;
  assign OptimizationBarrier_20_sum = TLB_covSum + OptimizationBarrier_20_io_covSum;
  assign OptimizationBarrier_21_sum = OptimizationBarrier_20_sum + OptimizationBarrier_21_io_covSum;
  assign OptimizationBarrier_35_sum = OptimizationBarrier_21_sum + OptimizationBarrier_35_io_covSum;
  assign OptimizationBarrier_6_sum = OptimizationBarrier_35_sum + OptimizationBarrier_6_io_covSum;
  assign OptimizationBarrier_16_sum = OptimizationBarrier_6_sum + OptimizationBarrier_16_io_covSum;
  assign OptimizationBarrier_12_sum = OptimizationBarrier_16_sum + OptimizationBarrier_12_io_covSum;
  assign OptimizationBarrier_9_sum = OptimizationBarrier_12_sum + OptimizationBarrier_9_io_covSum;
  assign OptimizationBarrier_8_sum = OptimizationBarrier_9_sum + OptimizationBarrier_8_io_covSum;
  assign OptimizationBarrier_2_sum = OptimizationBarrier_8_sum + OptimizationBarrier_2_io_covSum;
  assign OptimizationBarrier_25_sum = OptimizationBarrier_2_sum + OptimizationBarrier_25_io_covSum;
  assign pmp_sum = OptimizationBarrier_25_sum + pmp_io_covSum;
  assign OptimizationBarrier_23_sum = pmp_sum + OptimizationBarrier_23_io_covSum;
  assign OptimizationBarrier_27_sum = OptimizationBarrier_23_sum + OptimizationBarrier_27_io_covSum;
  assign OptimizationBarrier_30_sum = OptimizationBarrier_27_sum + OptimizationBarrier_30_io_covSum;
  assign OptimizationBarrier_1_sum = OptimizationBarrier_30_sum + OptimizationBarrier_1_io_covSum;
  assign OptimizationBarrier_18_sum = OptimizationBarrier_1_sum + OptimizationBarrier_18_io_covSum;
  assign OptimizationBarrier_31_sum = OptimizationBarrier_18_sum + OptimizationBarrier_31_io_covSum;
  assign OptimizationBarrier_19_sum = OptimizationBarrier_31_sum + OptimizationBarrier_19_io_covSum;
  assign OptimizationBarrier_37_sum = OptimizationBarrier_19_sum + OptimizationBarrier_37_io_covSum;
  assign OptimizationBarrier_28_sum = OptimizationBarrier_37_sum + OptimizationBarrier_28_io_covSum;
  assign OptimizationBarrier_33_sum = OptimizationBarrier_28_sum + OptimizationBarrier_33_io_covSum;
  assign OptimizationBarrier_4_sum = OptimizationBarrier_33_sum + OptimizationBarrier_4_io_covSum;
  assign OptimizationBarrier_38_sum = OptimizationBarrier_4_sum + OptimizationBarrier_38_io_covSum;
  assign OptimizationBarrier_sum = OptimizationBarrier_38_sum + OptimizationBarrier_io_covSum;
  assign OptimizationBarrier_34_sum = OptimizationBarrier_sum + OptimizationBarrier_34_io_covSum;
  assign OptimizationBarrier_24_sum = OptimizationBarrier_34_sum + OptimizationBarrier_24_io_covSum;
  assign OptimizationBarrier_22_sum = OptimizationBarrier_24_sum + OptimizationBarrier_22_io_covSum;
  assign OptimizationBarrier_10_sum = OptimizationBarrier_22_sum + OptimizationBarrier_10_io_covSum;
  assign OptimizationBarrier_3_sum = OptimizationBarrier_10_sum + OptimizationBarrier_3_io_covSum;
  assign OptimizationBarrier_5_sum = OptimizationBarrier_3_sum + OptimizationBarrier_5_io_covSum;
  assign OptimizationBarrier_36_sum = OptimizationBarrier_5_sum + OptimizationBarrier_36_io_covSum;
  assign OptimizationBarrier_17_sum = OptimizationBarrier_36_sum + OptimizationBarrier_17_io_covSum;
  assign OptimizationBarrier_15_sum = OptimizationBarrier_17_sum + OptimizationBarrier_15_io_covSum;
  assign OptimizationBarrier_29_sum = OptimizationBarrier_15_sum + OptimizationBarrier_29_io_covSum;
  assign OptimizationBarrier_32_sum = OptimizationBarrier_29_sum + OptimizationBarrier_32_io_covSum;
  assign OptimizationBarrier_7_sum = OptimizationBarrier_32_sum + OptimizationBarrier_7_io_covSum;
  assign OptimizationBarrier_14_sum = OptimizationBarrier_7_sum + OptimizationBarrier_14_io_covSum;
  assign OptimizationBarrier_26_sum = OptimizationBarrier_14_sum + OptimizationBarrier_26_io_covSum;
  assign OptimizationBarrier_11_sum = OptimizationBarrier_26_sum + OptimizationBarrier_11_io_covSum;
  assign OptimizationBarrier_13_sum = OptimizationBarrier_11_sum + OptimizationBarrier_13_io_covSum;
  assign io_covSum = OptimizationBarrier_13_sum;
  assign stopEn0 = io_sfence_valid & ~_T_2454;
  assign OptimizationBarrier_38_metaAssert_wire = OptimizationBarrier_38_metaAssert;
  assign OptimizationBarrier_2_metaAssert_wire = OptimizationBarrier_2_metaAssert;
  assign OptimizationBarrier_26_metaAssert_wire = OptimizationBarrier_26_metaAssert;
  assign OptimizationBarrier_metaAssert_wire = OptimizationBarrier_metaAssert;
  assign OptimizationBarrier_7_metaAssert_wire = OptimizationBarrier_7_metaAssert;
  assign OptimizationBarrier_37_metaAssert_wire = OptimizationBarrier_37_metaAssert;
  assign OptimizationBarrier_24_metaAssert_wire = OptimizationBarrier_24_metaAssert;
  assign OptimizationBarrier_17_metaAssert_wire = OptimizationBarrier_17_metaAssert;
  assign OptimizationBarrier_34_metaAssert_wire = OptimizationBarrier_34_metaAssert;
  assign OptimizationBarrier_21_metaAssert_wire = OptimizationBarrier_21_metaAssert;
  assign OptimizationBarrier_28_metaAssert_wire = OptimizationBarrier_28_metaAssert;
  assign OptimizationBarrier_16_metaAssert_wire = OptimizationBarrier_16_metaAssert;
  assign OptimizationBarrier_5_metaAssert_wire = OptimizationBarrier_5_metaAssert;
  assign OptimizationBarrier_8_metaAssert_wire = OptimizationBarrier_8_metaAssert;
  assign OptimizationBarrier_1_metaAssert_wire = OptimizationBarrier_1_metaAssert;
  assign OptimizationBarrier_4_metaAssert_wire = OptimizationBarrier_4_metaAssert;
  assign OptimizationBarrier_33_metaAssert_wire = OptimizationBarrier_33_metaAssert;
  assign OptimizationBarrier_30_metaAssert_wire = OptimizationBarrier_30_metaAssert;
  assign OptimizationBarrier_19_metaAssert_wire = OptimizationBarrier_19_metaAssert;
  assign OptimizationBarrier_20_metaAssert_wire = OptimizationBarrier_20_metaAssert;
  assign OptimizationBarrier_9_metaAssert_wire = OptimizationBarrier_9_metaAssert;
  assign OptimizationBarrier_29_metaAssert_wire = OptimizationBarrier_29_metaAssert;
  assign OptimizationBarrier_36_metaAssert_wire = OptimizationBarrier_36_metaAssert;
  assign OptimizationBarrier_31_metaAssert_wire = OptimizationBarrier_31_metaAssert;
  assign OptimizationBarrier_18_metaAssert_wire = OptimizationBarrier_18_metaAssert;
  assign OptimizationBarrier_12_metaAssert_wire = OptimizationBarrier_12_metaAssert;
  assign OptimizationBarrier_23_metaAssert_wire = OptimizationBarrier_23_metaAssert;
  assign OptimizationBarrier_32_metaAssert_wire = OptimizationBarrier_32_metaAssert;
  assign OptimizationBarrier_25_metaAssert_wire = OptimizationBarrier_25_metaAssert;
  assign pmp_metaAssert_wire = pmp_metaAssert;
  assign OptimizationBarrier_6_metaAssert_wire = OptimizationBarrier_6_metaAssert;
  assign OptimizationBarrier_27_metaAssert_wire = OptimizationBarrier_27_metaAssert;
  assign OptimizationBarrier_3_metaAssert_wire = OptimizationBarrier_3_metaAssert;
  assign OptimizationBarrier_14_metaAssert_wire = OptimizationBarrier_14_metaAssert;
  assign OptimizationBarrier_11_metaAssert_wire = OptimizationBarrier_11_metaAssert;
  assign OptimizationBarrier_15_metaAssert_wire = OptimizationBarrier_15_metaAssert;
  assign OptimizationBarrier_13_metaAssert_wire = OptimizationBarrier_13_metaAssert;
  assign OptimizationBarrier_22_metaAssert_wire = OptimizationBarrier_22_metaAssert;
  assign OptimizationBarrier_35_metaAssert_wire = OptimizationBarrier_35_metaAssert;
  assign OptimizationBarrier_10_metaAssert_wire = OptimizationBarrier_10_metaAssert;
  assign TLB_or15 = stopEn0 | OptimizationBarrier_33_metaAssert_wire;
  assign TLB_or34 = OptimizationBarrier_5_metaAssert_wire | OptimizationBarrier_20_metaAssert_wire;
  assign TLB_or16 = OptimizationBarrier_7_metaAssert_wire | TLB_or34;
  assign TLB_or7 = TLB_or15 | TLB_or16;
  assign TLB_or17 = OptimizationBarrier_22_metaAssert_wire | OptimizationBarrier_14_metaAssert_wire;
  assign TLB_or38 = OptimizationBarrier_metaAssert_wire | OptimizationBarrier_31_metaAssert_wire;
  assign TLB_or18 = OptimizationBarrier_2_metaAssert_wire | TLB_or38;
  assign TLB_or8 = TLB_or17 | TLB_or18;
  assign TLB_or3 = TLB_or7 | TLB_or8;
  assign TLB_or19 = OptimizationBarrier_18_metaAssert_wire | OptimizationBarrier_24_metaAssert_wire;
  assign TLB_or42 = OptimizationBarrier_25_metaAssert_wire | OptimizationBarrier_13_metaAssert_wire;
  assign TLB_or20 = OptimizationBarrier_10_metaAssert_wire | TLB_or42;
  assign TLB_or9 = TLB_or19 | TLB_or20;
  assign TLB_or21 = OptimizationBarrier_36_metaAssert_wire | OptimizationBarrier_34_metaAssert_wire;
  assign TLB_or46 = OptimizationBarrier_8_metaAssert_wire | OptimizationBarrier_21_metaAssert_wire;
  assign TLB_or22 = OptimizationBarrier_16_metaAssert_wire | TLB_or46;
  assign TLB_or10 = TLB_or21 | TLB_or22;
  assign TLB_or4 = TLB_or9 | TLB_or10;
  assign TLB_or1 = TLB_or3 | TLB_or4;
  assign TLB_or23 = OptimizationBarrier_12_metaAssert_wire | OptimizationBarrier_30_metaAssert_wire;
  assign TLB_or50 = OptimizationBarrier_27_metaAssert_wire | OptimizationBarrier_32_metaAssert_wire;
  assign TLB_or24 = pmp_metaAssert_wire | TLB_or50;
  assign TLB_or11 = TLB_or23 | TLB_or24;
  assign TLB_or25 = OptimizationBarrier_29_metaAssert_wire | OptimizationBarrier_1_metaAssert_wire;
  assign TLB_or54 = OptimizationBarrier_3_metaAssert_wire | OptimizationBarrier_38_metaAssert_wire;
  assign TLB_or26 = OptimizationBarrier_9_metaAssert_wire | TLB_or54;
  assign TLB_or12 = TLB_or25 | TLB_or26;
  assign TLB_or5 = TLB_or11 | TLB_or12;
  assign TLB_or27 = OptimizationBarrier_4_metaAssert_wire | OptimizationBarrier_6_metaAssert_wire;
  assign TLB_or58 = OptimizationBarrier_26_metaAssert_wire | OptimizationBarrier_19_metaAssert_wire;
  assign TLB_or28 = OptimizationBarrier_37_metaAssert_wire | TLB_or58;
  assign TLB_or13 = TLB_or27 | TLB_or28;
  assign TLB_or60 = OptimizationBarrier_11_metaAssert_wire | OptimizationBarrier_15_metaAssert_wire;
  assign TLB_or29 = OptimizationBarrier_28_metaAssert_wire | TLB_or60;
  assign TLB_or62 = OptimizationBarrier_17_metaAssert_wire | OptimizationBarrier_35_metaAssert_wire;
  assign TLB_or30 = OptimizationBarrier_23_metaAssert_wire | TLB_or62;
  assign TLB_or14 = TLB_or29 | TLB_or30;
  assign TLB_or6 = TLB_or13 | TLB_or14;
  assign TLB_or2 = TLB_or5 | TLB_or6;
  assign TLB_or0 = TLB_or1 | TLB_or2;
  assign metaAssert = TLB_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_tag = _RAND_0[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_data_0 = _RAND_1[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_data_1 = _RAND_2[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_data_2 = _RAND_3[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_data_3 = _RAND_4[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_valid_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_valid_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_valid_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_valid_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_1_tag = _RAND_9[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_1_data_0 = _RAND_10[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_1_data_1 = _RAND_11[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_1_data_2 = _RAND_12[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_1_data_3 = _RAND_13[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_1_valid_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_1_valid_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_1_valid_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_1_valid_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sectored_entries_2_tag = _RAND_18[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  sectored_entries_2_data_0 = _RAND_19[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  sectored_entries_2_data_1 = _RAND_20[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  sectored_entries_2_data_2 = _RAND_21[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  sectored_entries_2_data_3 = _RAND_22[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sectored_entries_2_valid_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sectored_entries_2_valid_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sectored_entries_2_valid_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sectored_entries_2_valid_3 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sectored_entries_3_tag = _RAND_27[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  sectored_entries_3_data_0 = _RAND_28[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  sectored_entries_3_data_1 = _RAND_29[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  sectored_entries_3_data_2 = _RAND_30[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  sectored_entries_3_data_3 = _RAND_31[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sectored_entries_3_valid_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sectored_entries_3_valid_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  sectored_entries_3_valid_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  sectored_entries_3_valid_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sectored_entries_4_tag = _RAND_36[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  sectored_entries_4_data_0 = _RAND_37[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  sectored_entries_4_data_1 = _RAND_38[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  sectored_entries_4_data_2 = _RAND_39[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  sectored_entries_4_data_3 = _RAND_40[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  sectored_entries_4_valid_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  sectored_entries_4_valid_1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  sectored_entries_4_valid_2 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  sectored_entries_4_valid_3 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  sectored_entries_5_tag = _RAND_45[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  sectored_entries_5_data_0 = _RAND_46[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  sectored_entries_5_data_1 = _RAND_47[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  sectored_entries_5_data_2 = _RAND_48[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  sectored_entries_5_data_3 = _RAND_49[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  sectored_entries_5_valid_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  sectored_entries_5_valid_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  sectored_entries_5_valid_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  sectored_entries_5_valid_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  sectored_entries_6_tag = _RAND_54[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  sectored_entries_6_data_0 = _RAND_55[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  sectored_entries_6_data_1 = _RAND_56[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  sectored_entries_6_data_2 = _RAND_57[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  sectored_entries_6_data_3 = _RAND_58[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  sectored_entries_6_valid_0 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  sectored_entries_6_valid_1 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  sectored_entries_6_valid_2 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  sectored_entries_6_valid_3 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  sectored_entries_7_tag = _RAND_63[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{`RANDOM}};
  sectored_entries_7_data_0 = _RAND_64[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  sectored_entries_7_data_1 = _RAND_65[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  sectored_entries_7_data_2 = _RAND_66[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  sectored_entries_7_data_3 = _RAND_67[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  sectored_entries_7_valid_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  sectored_entries_7_valid_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  sectored_entries_7_valid_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  sectored_entries_7_valid_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  superpage_entries_0_level = _RAND_72[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_73[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_74[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  superpage_entries_1_level = _RAND_76[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_77[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_78[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  superpage_entries_2_level = _RAND_80[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_81[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_82[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  superpage_entries_3_level = _RAND_84[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_85[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_86[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  special_entry_level = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  special_entry_tag = _RAND_89[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_90[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  state = _RAND_92[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  r_refill_tag = _RAND_93[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_94[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_96[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  r_sectored_hit = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_2116 = _RAND_98[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_2117 = _RAND_99[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  TLB_state = _RAND_100[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    TLB_cov[initvar] = _RAND_101[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  TLB_covSum = _RAND_102[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  TLB_metaAssert = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      sectored_entries_0_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1147) begin
            sectored_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1147) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1147) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1147) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1147) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2462) begin
          if (sectored_entries_0_data_0[0]) begin
            sectored_entries_0_valid_0 <= 1'h0;
          end else if (_T_422) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_0_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1147) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_valid_0 <= _GEN_85;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_0 <= _GEN_85;
                  end
                end
              end
            end
          end
        end else if (_T_422) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_0_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_0 <= _GEN_85;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1147) begin
                if (invalidate_refill) begin
                  sectored_entries_0_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_valid_0 <= _GEN_85;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_0 <= _GEN_685;
      end
    end else begin
      sectored_entries_0_valid_0 <= _GEN_505;
    end
    if (metaReset) begin
      sectored_entries_0_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_0_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2462) begin
          if (sectored_entries_0_data_1[0]) begin
            sectored_entries_0_valid_1 <= 1'h0;
          end else if (_T_422) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_0_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1147) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_valid_1 <= _GEN_86;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_1 <= _GEN_86;
                  end
                end
              end
            end
          end
        end else if (_T_422) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_0_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_1 <= _GEN_86;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1147) begin
                if (invalidate_refill) begin
                  sectored_entries_0_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_valid_1 <= _GEN_86;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_1 <= _GEN_686;
      end
    end else begin
      sectored_entries_0_valid_1 <= _GEN_506;
    end
    if (metaReset) begin
      sectored_entries_0_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_0_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2462) begin
          if (sectored_entries_0_data_2[0]) begin
            sectored_entries_0_valid_2 <= 1'h0;
          end else if (_T_422) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_0_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1147) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_valid_2 <= _GEN_87;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_2 <= _GEN_87;
                  end
                end
              end
            end
          end
        end else if (_T_422) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_0_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_2 <= _GEN_87;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1147) begin
                if (invalidate_refill) begin
                  sectored_entries_0_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_valid_2 <= _GEN_87;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_2 <= _GEN_687;
      end
    end else begin
      sectored_entries_0_valid_2 <= _GEN_507;
    end
    if (metaReset) begin
      sectored_entries_0_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_0_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2462) begin
          if (sectored_entries_0_data_3[0]) begin
            sectored_entries_0_valid_3 <= 1'h0;
          end else if (_T_422) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_0_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1147) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_valid_3 <= _GEN_88;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_3 <= _GEN_88;
                  end
                end
              end
            end
          end
        end else if (_T_422) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_0_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_3 <= _GEN_88;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1147) begin
                if (invalidate_refill) begin
                  sectored_entries_0_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_valid_3 <= _GEN_88;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_3 <= _GEN_688;
      end
    end else begin
      sectored_entries_0_valid_3 <= _GEN_508;
    end
    if (metaReset) begin
      sectored_entries_1_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1165) begin
            sectored_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1165) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1165) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1165) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1165) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2617) begin
          if (sectored_entries_1_data_0[0]) begin
            sectored_entries_1_valid_0 <= 1'h0;
          end else if (_T_428) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_1_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1165) begin
                    if (invalidate_refill) begin
                      sectored_entries_1_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_1_valid_0 <= _GEN_111;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_0 <= _GEN_111;
                  end
                end
              end
            end
          end
        end else if (_T_428) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_1_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_0 <= _GEN_111;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1165) begin
                if (invalidate_refill) begin
                  sectored_entries_1_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_1_valid_0 <= _GEN_111;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_0 <= _GEN_713;
      end
    end else begin
      sectored_entries_1_valid_0 <= _GEN_515;
    end
    if (metaReset) begin
      sectored_entries_1_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_1_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2617) begin
          if (sectored_entries_1_data_1[0]) begin
            sectored_entries_1_valid_1 <= 1'h0;
          end else if (_T_428) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_1_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1165) begin
                    if (invalidate_refill) begin
                      sectored_entries_1_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_1_valid_1 <= _GEN_112;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_1 <= _GEN_112;
                  end
                end
              end
            end
          end
        end else if (_T_428) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_1_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_1 <= _GEN_112;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1165) begin
                if (invalidate_refill) begin
                  sectored_entries_1_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_1_valid_1 <= _GEN_112;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_1 <= _GEN_714;
      end
    end else begin
      sectored_entries_1_valid_1 <= _GEN_516;
    end
    if (metaReset) begin
      sectored_entries_1_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_1_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2617) begin
          if (sectored_entries_1_data_2[0]) begin
            sectored_entries_1_valid_2 <= 1'h0;
          end else if (_T_428) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_1_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1165) begin
                    if (invalidate_refill) begin
                      sectored_entries_1_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_1_valid_2 <= _GEN_113;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_2 <= _GEN_113;
                  end
                end
              end
            end
          end
        end else if (_T_428) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_1_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_2 <= _GEN_113;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1165) begin
                if (invalidate_refill) begin
                  sectored_entries_1_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_1_valid_2 <= _GEN_113;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_2 <= _GEN_715;
      end
    end else begin
      sectored_entries_1_valid_2 <= _GEN_517;
    end
    if (metaReset) begin
      sectored_entries_1_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_1_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2617) begin
          if (sectored_entries_1_data_3[0]) begin
            sectored_entries_1_valid_3 <= 1'h0;
          end else if (_T_428) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_1_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1165) begin
                    if (invalidate_refill) begin
                      sectored_entries_1_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_1_valid_3 <= _GEN_114;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_3 <= _GEN_114;
                  end
                end
              end
            end
          end
        end else if (_T_428) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_1_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_3 <= _GEN_114;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1165) begin
                if (invalidate_refill) begin
                  sectored_entries_1_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_1_valid_3 <= _GEN_114;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_3 <= _GEN_716;
      end
    end else begin
      sectored_entries_1_valid_3 <= _GEN_518;
    end
    if (metaReset) begin
      sectored_entries_2_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1183) begin
            sectored_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1183) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1183) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1183) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1183) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2772) begin
          if (sectored_entries_2_data_0[0]) begin
            sectored_entries_2_valid_0 <= 1'h0;
          end else if (_T_434) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_2_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1183) begin
                    if (invalidate_refill) begin
                      sectored_entries_2_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_2_valid_0 <= _GEN_137;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_0 <= _GEN_137;
                  end
                end
              end
            end
          end
        end else if (_T_434) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_2_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_0 <= _GEN_137;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1183) begin
                if (invalidate_refill) begin
                  sectored_entries_2_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_2_valid_0 <= _GEN_137;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_0 <= _GEN_741;
      end
    end else begin
      sectored_entries_2_valid_0 <= _GEN_525;
    end
    if (metaReset) begin
      sectored_entries_2_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_2_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2772) begin
          if (sectored_entries_2_data_1[0]) begin
            sectored_entries_2_valid_1 <= 1'h0;
          end else if (_T_434) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_2_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1183) begin
                    if (invalidate_refill) begin
                      sectored_entries_2_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_2_valid_1 <= _GEN_138;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_1 <= _GEN_138;
                  end
                end
              end
            end
          end
        end else if (_T_434) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_2_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_1 <= _GEN_138;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1183) begin
                if (invalidate_refill) begin
                  sectored_entries_2_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_2_valid_1 <= _GEN_138;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_1 <= _GEN_742;
      end
    end else begin
      sectored_entries_2_valid_1 <= _GEN_526;
    end
    if (metaReset) begin
      sectored_entries_2_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_2_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2772) begin
          if (sectored_entries_2_data_2[0]) begin
            sectored_entries_2_valid_2 <= 1'h0;
          end else if (_T_434) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_2_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1183) begin
                    if (invalidate_refill) begin
                      sectored_entries_2_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_2_valid_2 <= _GEN_139;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_2 <= _GEN_139;
                  end
                end
              end
            end
          end
        end else if (_T_434) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_2_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_2 <= _GEN_139;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1183) begin
                if (invalidate_refill) begin
                  sectored_entries_2_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_2_valid_2 <= _GEN_139;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_2 <= _GEN_743;
      end
    end else begin
      sectored_entries_2_valid_2 <= _GEN_527;
    end
    if (metaReset) begin
      sectored_entries_2_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_2_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2772) begin
          if (sectored_entries_2_data_3[0]) begin
            sectored_entries_2_valid_3 <= 1'h0;
          end else if (_T_434) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_2_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1183) begin
                    if (invalidate_refill) begin
                      sectored_entries_2_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_2_valid_3 <= _GEN_140;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_3 <= _GEN_140;
                  end
                end
              end
            end
          end
        end else if (_T_434) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_2_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_3 <= _GEN_140;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1183) begin
                if (invalidate_refill) begin
                  sectored_entries_2_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_2_valid_3 <= _GEN_140;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_3 <= _GEN_744;
      end
    end else begin
      sectored_entries_2_valid_3 <= _GEN_528;
    end
    if (metaReset) begin
      sectored_entries_3_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1201) begin
            sectored_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1201) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1201) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1201) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1201) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2927) begin
          if (sectored_entries_3_data_0[0]) begin
            sectored_entries_3_valid_0 <= 1'h0;
          end else if (_T_440) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_3_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1201) begin
                    if (invalidate_refill) begin
                      sectored_entries_3_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_3_valid_0 <= _GEN_163;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_0 <= _GEN_163;
                  end
                end
              end
            end
          end
        end else if (_T_440) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_3_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_0 <= _GEN_163;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1201) begin
                if (invalidate_refill) begin
                  sectored_entries_3_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_3_valid_0 <= _GEN_163;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_0 <= _GEN_769;
      end
    end else begin
      sectored_entries_3_valid_0 <= _GEN_535;
    end
    if (metaReset) begin
      sectored_entries_3_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_3_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2927) begin
          if (sectored_entries_3_data_1[0]) begin
            sectored_entries_3_valid_1 <= 1'h0;
          end else if (_T_440) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_3_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1201) begin
                    if (invalidate_refill) begin
                      sectored_entries_3_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_3_valid_1 <= _GEN_164;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_1 <= _GEN_164;
                  end
                end
              end
            end
          end
        end else if (_T_440) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_3_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_1 <= _GEN_164;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1201) begin
                if (invalidate_refill) begin
                  sectored_entries_3_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_3_valid_1 <= _GEN_164;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_1 <= _GEN_770;
      end
    end else begin
      sectored_entries_3_valid_1 <= _GEN_536;
    end
    if (metaReset) begin
      sectored_entries_3_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_3_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2927) begin
          if (sectored_entries_3_data_2[0]) begin
            sectored_entries_3_valid_2 <= 1'h0;
          end else if (_T_440) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_3_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1201) begin
                    if (invalidate_refill) begin
                      sectored_entries_3_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_3_valid_2 <= _GEN_165;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_2 <= _GEN_165;
                  end
                end
              end
            end
          end
        end else if (_T_440) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_3_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_2 <= _GEN_165;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1201) begin
                if (invalidate_refill) begin
                  sectored_entries_3_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_3_valid_2 <= _GEN_165;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_2 <= _GEN_771;
      end
    end else begin
      sectored_entries_3_valid_2 <= _GEN_537;
    end
    if (metaReset) begin
      sectored_entries_3_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_3_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2927) begin
          if (sectored_entries_3_data_3[0]) begin
            sectored_entries_3_valid_3 <= 1'h0;
          end else if (_T_440) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_3_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1201) begin
                    if (invalidate_refill) begin
                      sectored_entries_3_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_3_valid_3 <= _GEN_166;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_3 <= _GEN_166;
                  end
                end
              end
            end
          end
        end else if (_T_440) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_3_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_3 <= _GEN_166;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1201) begin
                if (invalidate_refill) begin
                  sectored_entries_3_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_3_valid_3 <= _GEN_166;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_3 <= _GEN_772;
      end
    end else begin
      sectored_entries_3_valid_3 <= _GEN_538;
    end
    if (metaReset) begin
      sectored_entries_4_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1219) begin
            sectored_entries_4_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1219) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1219) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1219) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1219) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_4_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3082) begin
          if (sectored_entries_4_data_0[0]) begin
            sectored_entries_4_valid_0 <= 1'h0;
          end else if (_T_446) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_4_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1219) begin
                    if (invalidate_refill) begin
                      sectored_entries_4_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_4_valid_0 <= _GEN_189;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_0 <= _GEN_189;
                  end
                end
              end
            end
          end
        end else if (_T_446) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_4_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_0 <= _GEN_189;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1219) begin
                if (invalidate_refill) begin
                  sectored_entries_4_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_4_valid_0 <= _GEN_189;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_0 <= _GEN_797;
      end
    end else begin
      sectored_entries_4_valid_0 <= _GEN_545;
    end
    if (metaReset) begin
      sectored_entries_4_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_4_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3082) begin
          if (sectored_entries_4_data_1[0]) begin
            sectored_entries_4_valid_1 <= 1'h0;
          end else if (_T_446) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_4_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1219) begin
                    if (invalidate_refill) begin
                      sectored_entries_4_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_4_valid_1 <= _GEN_190;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_1 <= _GEN_190;
                  end
                end
              end
            end
          end
        end else if (_T_446) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_4_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_1 <= _GEN_190;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1219) begin
                if (invalidate_refill) begin
                  sectored_entries_4_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_4_valid_1 <= _GEN_190;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_1 <= _GEN_798;
      end
    end else begin
      sectored_entries_4_valid_1 <= _GEN_546;
    end
    if (metaReset) begin
      sectored_entries_4_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_4_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3082) begin
          if (sectored_entries_4_data_2[0]) begin
            sectored_entries_4_valid_2 <= 1'h0;
          end else if (_T_446) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_4_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1219) begin
                    if (invalidate_refill) begin
                      sectored_entries_4_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_4_valid_2 <= _GEN_191;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_2 <= _GEN_191;
                  end
                end
              end
            end
          end
        end else if (_T_446) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_4_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_2 <= _GEN_191;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1219) begin
                if (invalidate_refill) begin
                  sectored_entries_4_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_4_valid_2 <= _GEN_191;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_2 <= _GEN_799;
      end
    end else begin
      sectored_entries_4_valid_2 <= _GEN_547;
    end
    if (metaReset) begin
      sectored_entries_4_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_4_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3082) begin
          if (sectored_entries_4_data_3[0]) begin
            sectored_entries_4_valid_3 <= 1'h0;
          end else if (_T_446) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_4_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1219) begin
                    if (invalidate_refill) begin
                      sectored_entries_4_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_4_valid_3 <= _GEN_192;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_3 <= _GEN_192;
                  end
                end
              end
            end
          end
        end else if (_T_446) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_4_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_3 <= _GEN_192;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1219) begin
                if (invalidate_refill) begin
                  sectored_entries_4_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_4_valid_3 <= _GEN_192;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_3 <= _GEN_800;
      end
    end else begin
      sectored_entries_4_valid_3 <= _GEN_548;
    end
    if (metaReset) begin
      sectored_entries_5_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1237) begin
            sectored_entries_5_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1237) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1237) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1237) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1237) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_5_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3237) begin
          if (sectored_entries_5_data_0[0]) begin
            sectored_entries_5_valid_0 <= 1'h0;
          end else if (_T_452) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_5_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1237) begin
                    if (invalidate_refill) begin
                      sectored_entries_5_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_5_valid_0 <= _GEN_215;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_0 <= _GEN_215;
                  end
                end
              end
            end
          end
        end else if (_T_452) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_5_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_0 <= _GEN_215;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1237) begin
                if (invalidate_refill) begin
                  sectored_entries_5_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_5_valid_0 <= _GEN_215;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_0 <= _GEN_825;
      end
    end else begin
      sectored_entries_5_valid_0 <= _GEN_555;
    end
    if (metaReset) begin
      sectored_entries_5_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_5_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3237) begin
          if (sectored_entries_5_data_1[0]) begin
            sectored_entries_5_valid_1 <= 1'h0;
          end else if (_T_452) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_5_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1237) begin
                    if (invalidate_refill) begin
                      sectored_entries_5_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_5_valid_1 <= _GEN_216;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_1 <= _GEN_216;
                  end
                end
              end
            end
          end
        end else if (_T_452) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_5_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_1 <= _GEN_216;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1237) begin
                if (invalidate_refill) begin
                  sectored_entries_5_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_5_valid_1 <= _GEN_216;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_1 <= _GEN_826;
      end
    end else begin
      sectored_entries_5_valid_1 <= _GEN_556;
    end
    if (metaReset) begin
      sectored_entries_5_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_5_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3237) begin
          if (sectored_entries_5_data_2[0]) begin
            sectored_entries_5_valid_2 <= 1'h0;
          end else if (_T_452) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_5_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1237) begin
                    if (invalidate_refill) begin
                      sectored_entries_5_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_5_valid_2 <= _GEN_217;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_2 <= _GEN_217;
                  end
                end
              end
            end
          end
        end else if (_T_452) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_5_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_2 <= _GEN_217;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1237) begin
                if (invalidate_refill) begin
                  sectored_entries_5_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_5_valid_2 <= _GEN_217;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_2 <= _GEN_827;
      end
    end else begin
      sectored_entries_5_valid_2 <= _GEN_557;
    end
    if (metaReset) begin
      sectored_entries_5_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_5_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3237) begin
          if (sectored_entries_5_data_3[0]) begin
            sectored_entries_5_valid_3 <= 1'h0;
          end else if (_T_452) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_5_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1237) begin
                    if (invalidate_refill) begin
                      sectored_entries_5_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_5_valid_3 <= _GEN_218;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_3 <= _GEN_218;
                  end
                end
              end
            end
          end
        end else if (_T_452) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_5_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_3 <= _GEN_218;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1237) begin
                if (invalidate_refill) begin
                  sectored_entries_5_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_5_valid_3 <= _GEN_218;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_3 <= _GEN_828;
      end
    end else begin
      sectored_entries_5_valid_3 <= _GEN_558;
    end
    if (metaReset) begin
      sectored_entries_6_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1255) begin
            sectored_entries_6_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1255) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1255) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1255) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1255) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_6_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3392) begin
          if (sectored_entries_6_data_0[0]) begin
            sectored_entries_6_valid_0 <= 1'h0;
          end else if (_T_458) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_6_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1255) begin
                    if (invalidate_refill) begin
                      sectored_entries_6_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_6_valid_0 <= _GEN_241;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_0 <= _GEN_241;
                  end
                end
              end
            end
          end
        end else if (_T_458) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_6_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_0 <= _GEN_241;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1255) begin
                if (invalidate_refill) begin
                  sectored_entries_6_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_6_valid_0 <= _GEN_241;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_0 <= _GEN_853;
      end
    end else begin
      sectored_entries_6_valid_0 <= _GEN_565;
    end
    if (metaReset) begin
      sectored_entries_6_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_6_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3392) begin
          if (sectored_entries_6_data_1[0]) begin
            sectored_entries_6_valid_1 <= 1'h0;
          end else if (_T_458) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_6_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1255) begin
                    if (invalidate_refill) begin
                      sectored_entries_6_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_6_valid_1 <= _GEN_242;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_1 <= _GEN_242;
                  end
                end
              end
            end
          end
        end else if (_T_458) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_6_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_1 <= _GEN_242;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1255) begin
                if (invalidate_refill) begin
                  sectored_entries_6_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_6_valid_1 <= _GEN_242;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_1 <= _GEN_854;
      end
    end else begin
      sectored_entries_6_valid_1 <= _GEN_566;
    end
    if (metaReset) begin
      sectored_entries_6_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_6_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3392) begin
          if (sectored_entries_6_data_2[0]) begin
            sectored_entries_6_valid_2 <= 1'h0;
          end else if (_T_458) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_6_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1255) begin
                    if (invalidate_refill) begin
                      sectored_entries_6_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_6_valid_2 <= _GEN_243;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_2 <= _GEN_243;
                  end
                end
              end
            end
          end
        end else if (_T_458) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_6_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_2 <= _GEN_243;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1255) begin
                if (invalidate_refill) begin
                  sectored_entries_6_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_6_valid_2 <= _GEN_243;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_2 <= _GEN_855;
      end
    end else begin
      sectored_entries_6_valid_2 <= _GEN_567;
    end
    if (metaReset) begin
      sectored_entries_6_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_6_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3392) begin
          if (sectored_entries_6_data_3[0]) begin
            sectored_entries_6_valid_3 <= 1'h0;
          end else if (_T_458) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_6_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1255) begin
                    if (invalidate_refill) begin
                      sectored_entries_6_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_6_valid_3 <= _GEN_244;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_3 <= _GEN_244;
                  end
                end
              end
            end
          end
        end else if (_T_458) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_6_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_3 <= _GEN_244;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1255) begin
                if (invalidate_refill) begin
                  sectored_entries_6_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_6_valid_3 <= _GEN_244;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_3 <= _GEN_856;
      end
    end else begin
      sectored_entries_6_valid_3 <= _GEN_568;
    end
    if (metaReset) begin
      sectored_entries_7_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1273) begin
            sectored_entries_7_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1273) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1273) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1273) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1273) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_7_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3547) begin
          if (sectored_entries_7_data_0[0]) begin
            sectored_entries_7_valid_0 <= 1'h0;
          end else if (_T_464) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_7_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1273) begin
                    if (invalidate_refill) begin
                      sectored_entries_7_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_7_valid_0 <= _GEN_267;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_0 <= _GEN_267;
                  end
                end
              end
            end
          end
        end else if (_T_464) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_7_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_0 <= _GEN_267;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1273) begin
                if (invalidate_refill) begin
                  sectored_entries_7_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_7_valid_0 <= _GEN_267;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_0 <= _GEN_881;
      end
    end else begin
      sectored_entries_7_valid_0 <= _GEN_575;
    end
    if (metaReset) begin
      sectored_entries_7_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_7_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3547) begin
          if (sectored_entries_7_data_1[0]) begin
            sectored_entries_7_valid_1 <= 1'h0;
          end else if (_T_464) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_7_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1273) begin
                    if (invalidate_refill) begin
                      sectored_entries_7_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_7_valid_1 <= _GEN_268;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_1 <= _GEN_268;
                  end
                end
              end
            end
          end
        end else if (_T_464) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_7_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_1 <= _GEN_268;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1273) begin
                if (invalidate_refill) begin
                  sectored_entries_7_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_7_valid_1 <= _GEN_268;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_1 <= _GEN_882;
      end
    end else begin
      sectored_entries_7_valid_1 <= _GEN_576;
    end
    if (metaReset) begin
      sectored_entries_7_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_7_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3547) begin
          if (sectored_entries_7_data_2[0]) begin
            sectored_entries_7_valid_2 <= 1'h0;
          end else if (_T_464) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_7_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1273) begin
                    if (invalidate_refill) begin
                      sectored_entries_7_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_7_valid_2 <= _GEN_269;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_2 <= _GEN_269;
                  end
                end
              end
            end
          end
        end else if (_T_464) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_7_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_2 <= _GEN_269;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1273) begin
                if (invalidate_refill) begin
                  sectored_entries_7_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_7_valid_2 <= _GEN_269;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_2 <= _GEN_883;
      end
    end else begin
      sectored_entries_7_valid_2 <= _GEN_577;
    end
    if (metaReset) begin
      sectored_entries_7_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_7_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3547) begin
          if (sectored_entries_7_data_3[0]) begin
            sectored_entries_7_valid_3 <= 1'h0;
          end else if (_T_464) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_7_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1273) begin
                    if (invalidate_refill) begin
                      sectored_entries_7_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_7_valid_3 <= _GEN_270;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_3 <= _GEN_270;
                  end
                end
              end
            end
          end
        end else if (_T_464) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_7_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_3 <= _GEN_270;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1273) begin
                if (invalidate_refill) begin
                  sectored_entries_7_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_7_valid_3 <= _GEN_270;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_3 <= _GEN_884;
      end
    end else begin
      sectored_entries_7_valid_3 <= _GEN_578;
    end
    if (metaReset) begin
      superpage_entries_0_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1078) begin
            superpage_entries_0_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1078) begin
            superpage_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1078) begin
            superpage_entries_0_data_0 <= _T_1076;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_0) begin
          superpage_entries_0_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1077) begin
              if (_T_1078) begin
                if (invalidate_refill) begin
                  superpage_entries_0_valid_0 <= 1'h0;
                end else begin
                  superpage_entries_0_valid_0 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        superpage_entries_0_valid_0 <= _GEN_891;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1078) begin
            if (invalidate_refill) begin
              superpage_entries_0_valid_0 <= 1'h0;
            end else begin
              superpage_entries_0_valid_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1095) begin
            superpage_entries_1_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1095) begin
            superpage_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1095) begin
            superpage_entries_1_data_0 <= _T_1076;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_1) begin
          superpage_entries_1_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1077) begin
              if (_T_1095) begin
                if (invalidate_refill) begin
                  superpage_entries_1_valid_0 <= 1'h0;
                end else begin
                  superpage_entries_1_valid_0 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        superpage_entries_1_valid_0 <= _GEN_895;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1095) begin
            if (invalidate_refill) begin
              superpage_entries_1_valid_0 <= 1'h0;
            end else begin
              superpage_entries_1_valid_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1112) begin
            superpage_entries_2_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1112) begin
            superpage_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1112) begin
            superpage_entries_2_data_0 <= _T_1076;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_2) begin
          superpage_entries_2_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1077) begin
              if (_T_1112) begin
                superpage_entries_2_valid_0 <= _GEN_64;
              end
            end
          end
        end
      end else begin
        superpage_entries_2_valid_0 <= _GEN_899;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1112) begin
            superpage_entries_2_valid_0 <= _GEN_64;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1129) begin
            superpage_entries_3_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1129) begin
            superpage_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1129) begin
            superpage_entries_3_data_0 <= _T_1076;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_3) begin
          superpage_entries_3_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1077) begin
              if (_T_1129) begin
                superpage_entries_3_valid_0 <= _GEN_64;
              end
            end
          end
        end
      end else begin
        superpage_entries_3_valid_0 <= _GEN_903;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1129) begin
            superpage_entries_3_valid_0 <= _GEN_64;
          end
        end
      end
    end
    if (metaReset) begin
      special_entry_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_level <= io_ptw_resp_bits_level;
      end
    end
    if (metaReset) begin
      special_entry_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_tag <= r_refill_tag;
      end
    end
    if (metaReset) begin
      special_entry_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_data_0 <= _T_1076;
      end
    end
    if (metaReset) begin
      special_entry_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      special_entry_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_689) begin
          special_entry_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (~io_ptw_resp_bits_homogeneous) begin
            special_entry_valid_0 <= _GEN_64;
          end
        end
      end else begin
        special_entry_valid_0 <= _GEN_907;
      end
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_valid_0 <= _GEN_64;
      end
    end
    if (metaReset) begin
      state <= 2'h0;
    end else if (reset) begin
      state <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if (_T_2448) begin
      state <= 2'h3;
    end else if (_T_4) begin
      if (io_ptw_req_ready) begin
        if (io_sfence_valid) begin
          state <= 2'h3;
        end else begin
          state <= 2'h2;
        end
      end else if (io_sfence_valid) begin
        state <= 2'h0;
      end else if (_T_2331) begin
        state <= 2'h1;
      end
    end else if (_T_2331) begin
      state <= 2'h1;
    end
    if (metaReset) begin
      r_refill_tag <= 27'h0;
    end else if (_T_2331) begin
      r_refill_tag <= vpn;
    end
    if (metaReset) begin
      r_superpage_repl_addr <= 2'h0;
    end else if (_T_2331) begin
      if (_T_2342) begin
        r_superpage_repl_addr <= _T_2338;
      end else if (_T_2344) begin
        r_superpage_repl_addr <= 2'h0;
      end else if (_T_2345) begin
        r_superpage_repl_addr <= 2'h1;
      end else if (_T_2346) begin
        r_superpage_repl_addr <= 2'h2;
      end else begin
        r_superpage_repl_addr <= 2'h3;
      end
    end
    if (metaReset) begin
      r_sectored_repl_addr <= 3'h0;
    end else if (_T_2331) begin
      if (_T_2402) begin
        r_sectored_repl_addr <= _T_2370;
      end else if (_T_2404) begin
        r_sectored_repl_addr <= 3'h0;
      end else if (_T_2405) begin
        r_sectored_repl_addr <= 3'h1;
      end else if (_T_2406) begin
        r_sectored_repl_addr <= 3'h2;
      end else if (_T_2407) begin
        r_sectored_repl_addr <= 3'h3;
      end else if (_T_2408) begin
        r_sectored_repl_addr <= 3'h4;
      end else if (_T_2409) begin
        r_sectored_repl_addr <= 3'h5;
      end else if (_T_2410) begin
        r_sectored_repl_addr <= 3'h6;
      end else begin
        r_sectored_repl_addr <= 3'h7;
      end
    end
    if (metaReset) begin
      r_sectored_hit_addr <= 3'h0;
    end else if (_T_2331) begin
      r_sectored_hit_addr <= _T_2143;
    end
    if (metaReset) begin
      r_sectored_hit <= 1'h0;
    end else if (_T_2331) begin
      r_sectored_hit <= _T_2125;
    end
    if (metaReset) begin
      _T_2116 <= 7'h0;
    end else if (_T_2118) begin
      if (_T_2125) begin
        _T_2116 <= _T_2182;
      end
    end
    if (metaReset) begin
      _T_2117 <= 3'h0;
    end else if (_T_2118) begin
      if (_T_2185) begin
        _T_2117 <= _T_2209;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & ~_T_2454) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:381 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"); // @[TLB.scala 381:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_sfence_valid & ~_T_2454) begin
          $fatal; // @[TLB.scala 381:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    TLB_state <= TLB_xor0;
    if (!(TLB_cov_read_data)) begin
      TLB_covSum <= TLB_covSum + 1'h1;
    end
    if (metaReset) begin
      TLB_metaAssert <= 1'h0;
    end else begin
      TLB_metaAssert <= TLB_metaAssert | TLB_or0;
    end
  end
  always @(posedge clock) begin
    if(TLB_cov_write_en & TLB_cov_write_mask) begin
      TLB_cov[TLB_cov_write_addr] <= TLB_cov_write_data; // @[Coverage map for TLB]
    end
  end
endmodule
module MaxPeriodFibonacciLFSR(
  input         clock,
  input         reset,
  input         io_increment,
  output        io_out_0,
  output        io_out_1,
  output        io_out_2,
  output        io_out_3,
  output        io_out_4,
  output        io_out_5,
  output        io_out_6,
  output        io_out_7,
  output        io_out_8,
  output        io_out_9,
  output        io_out_10,
  output        io_out_11,
  output        io_out_12,
  output        io_out_13,
  output        io_out_14,
  output        io_out_15,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  state_0; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_0;
  reg  state_1; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_1;
  reg  state_2; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_2;
  reg  state_3; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_3;
  reg  state_4; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_4;
  reg  state_5; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_5;
  reg  state_6; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_6;
  reg  state_7; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_7;
  reg  state_8; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_8;
  reg  state_9; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_9;
  reg  state_10; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_10;
  reg  state_11; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_11;
  reg  state_12; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_12;
  reg  state_13; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_13;
  reg  state_14; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_14;
  reg  state_15; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_15;
  wire  _T_1; // @[LFSR.scala 15:41]
  wire  _T_2; // @[LFSR.scala 15:41]
  wire  _T_3; // @[LFSR.scala 15:41]
  wire  _GEN_0; // @[PRNG.scala 61:23]
  wire [29:0] MaxPeriodFibonacciLFSR_covSum;
  assign _T_1 = state_15 ^ state_13; // @[LFSR.scala 15:41]
  assign _T_2 = _T_1 ^ state_12; // @[LFSR.scala 15:41]
  assign _T_3 = _T_2 ^ state_10; // @[LFSR.scala 15:41]
  assign _GEN_0 = io_increment ? _T_3 : state_0; // @[PRNG.scala 61:23]
  assign io_out_0 = state_0; // @[PRNG.scala 69:10]
  assign io_out_1 = state_1; // @[PRNG.scala 69:10]
  assign io_out_2 = state_2; // @[PRNG.scala 69:10]
  assign io_out_3 = state_3; // @[PRNG.scala 69:10]
  assign io_out_4 = state_4; // @[PRNG.scala 69:10]
  assign io_out_5 = state_5; // @[PRNG.scala 69:10]
  assign io_out_6 = state_6; // @[PRNG.scala 69:10]
  assign io_out_7 = state_7; // @[PRNG.scala 69:10]
  assign io_out_8 = state_8; // @[PRNG.scala 69:10]
  assign io_out_9 = state_9; // @[PRNG.scala 69:10]
  assign io_out_10 = state_10; // @[PRNG.scala 69:10]
  assign io_out_11 = state_11; // @[PRNG.scala 69:10]
  assign io_out_12 = state_12; // @[PRNG.scala 69:10]
  assign io_out_13 = state_13; // @[PRNG.scala 69:10]
  assign io_out_14 = state_14; // @[PRNG.scala 69:10]
  assign io_out_15 = state_15; // @[PRNG.scala 69:10]
  assign MaxPeriodFibonacciLFSR_covSum = 30'h0;
  assign io_covSum = MaxPeriodFibonacciLFSR_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      state_0 <= 1'h0;
    end else begin
      state_0 <= reset | _GEN_0;
    end
    if (metaReset) begin
      state_1 <= 1'h0;
    end else if (reset) begin
      state_1 <= 1'h0;
    end else if (io_increment) begin
      state_1 <= state_0;
    end
    if (metaReset) begin
      state_2 <= 1'h0;
    end else if (reset) begin
      state_2 <= 1'h0;
    end else if (io_increment) begin
      state_2 <= state_1;
    end
    if (metaReset) begin
      state_3 <= 1'h0;
    end else if (reset) begin
      state_3 <= 1'h0;
    end else if (io_increment) begin
      state_3 <= state_2;
    end
    if (metaReset) begin
      state_4 <= 1'h0;
    end else if (reset) begin
      state_4 <= 1'h0;
    end else if (io_increment) begin
      state_4 <= state_3;
    end
    if (metaReset) begin
      state_5 <= 1'h0;
    end else if (reset) begin
      state_5 <= 1'h0;
    end else if (io_increment) begin
      state_5 <= state_4;
    end
    if (metaReset) begin
      state_6 <= 1'h0;
    end else if (reset) begin
      state_6 <= 1'h0;
    end else if (io_increment) begin
      state_6 <= state_5;
    end
    if (metaReset) begin
      state_7 <= 1'h0;
    end else if (reset) begin
      state_7 <= 1'h0;
    end else if (io_increment) begin
      state_7 <= state_6;
    end
    if (metaReset) begin
      state_8 <= 1'h0;
    end else if (reset) begin
      state_8 <= 1'h0;
    end else if (io_increment) begin
      state_8 <= state_7;
    end
    if (metaReset) begin
      state_9 <= 1'h0;
    end else if (reset) begin
      state_9 <= 1'h0;
    end else if (io_increment) begin
      state_9 <= state_8;
    end
    if (metaReset) begin
      state_10 <= 1'h0;
    end else if (reset) begin
      state_10 <= 1'h0;
    end else if (io_increment) begin
      state_10 <= state_9;
    end
    if (metaReset) begin
      state_11 <= 1'h0;
    end else if (reset) begin
      state_11 <= 1'h0;
    end else if (io_increment) begin
      state_11 <= state_10;
    end
    if (metaReset) begin
      state_12 <= 1'h0;
    end else if (reset) begin
      state_12 <= 1'h0;
    end else if (io_increment) begin
      state_12 <= state_11;
    end
    if (metaReset) begin
      state_13 <= 1'h0;
    end else if (reset) begin
      state_13 <= 1'h0;
    end else if (io_increment) begin
      state_13 <= state_12;
    end
    if (metaReset) begin
      state_14 <= 1'h0;
    end else if (reset) begin
      state_14 <= 1'h0;
    end else if (io_increment) begin
      state_14 <= state_13;
    end
    if (metaReset) begin
      state_15 <= 1'h0;
    end else if (reset) begin
      state_15 <= 1'h0;
    end else if (io_increment) begin
      state_15 <= state_14;
    end
  end
endmodule
module DCacheModuleImpl_Anon_1(
  input         io_in_0_valid,
  input  [39:0] io_in_0_bits_addr,
  input  [5:0]  io_in_0_bits_idx,
  input  [21:0] io_in_0_bits_data,
  input         io_in_1_valid,
  input  [39:0] io_in_1_bits_addr,
  input  [5:0]  io_in_1_bits_idx,
  input  [21:0] io_in_1_bits_data,
  input         io_in_2_valid,
  input  [39:0] io_in_2_bits_addr,
  input  [5:0]  io_in_2_bits_idx,
  input  [3:0]  io_in_2_bits_way_en,
  input  [21:0] io_in_2_bits_data,
  input         io_in_3_valid,
  input  [39:0] io_in_3_bits_addr,
  input  [5:0]  io_in_3_bits_idx,
  input  [3:0]  io_in_3_bits_way_en,
  input  [21:0] io_in_3_bits_data,
  output        io_in_4_ready,
  input         io_in_4_valid,
  input  [39:0] io_in_4_bits_addr,
  input  [5:0]  io_in_4_bits_idx,
  input  [3:0]  io_in_4_bits_way_en,
  input  [21:0] io_in_4_bits_data,
  output        io_in_5_ready,
  input         io_in_5_valid,
  input  [39:0] io_in_5_bits_addr,
  input  [5:0]  io_in_5_bits_idx,
  output        io_in_6_ready,
  input         io_in_6_valid,
  input  [39:0] io_in_6_bits_addr,
  input  [5:0]  io_in_6_bits_idx,
  input  [3:0]  io_in_6_bits_way_en,
  input  [21:0] io_in_6_bits_data,
  output        io_in_7_ready,
  input         io_in_7_valid,
  input  [39:0] io_in_7_bits_addr,
  input  [5:0]  io_in_7_bits_idx,
  input  [3:0]  io_in_7_bits_way_en,
  input  [21:0] io_in_7_bits_data,
  output        io_out_valid,
  output        io_out_bits_write,
  output [39:0] io_out_bits_addr,
  output [5:0]  io_out_bits_idx,
  output [3:0]  io_out_bits_way_en,
  output [21:0] io_out_bits_data,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [21:0] _GEN_1; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_2; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_3; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_4; // @[Arbiter.scala 126:27]
  wire [21:0] _GEN_13; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_14; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_15; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_16; // @[Arbiter.scala 126:27]
  wire [21:0] _GEN_19; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_20; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_21; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_22; // @[Arbiter.scala 126:27]
  wire  _GEN_23; // @[Arbiter.scala 126:27]
  wire [21:0] _GEN_25; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_26; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_27; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_28; // @[Arbiter.scala 126:27]
  wire  _GEN_29; // @[Arbiter.scala 126:27]
  wire [21:0] _GEN_31; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_32; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_33; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_34; // @[Arbiter.scala 126:27]
  wire  _GEN_35; // @[Arbiter.scala 126:27]
  wire  _T; // @[Arbiter.scala 31:68]
  wire  _T_1; // @[Arbiter.scala 31:68]
  wire  _T_2; // @[Arbiter.scala 31:68]
  wire  _T_3; // @[Arbiter.scala 31:68]
  wire  _T_5; // @[Arbiter.scala 31:68]
  wire  grant_7; // @[Arbiter.scala 31:78]
  wire [29:0] DCacheModuleImpl_Anon_1_covSum;
  assign _GEN_1 = io_in_6_valid ? io_in_6_bits_data : io_in_7_bits_data; // @[Arbiter.scala 126:27]
  assign _GEN_2 = io_in_6_valid ? io_in_6_bits_way_en : io_in_7_bits_way_en; // @[Arbiter.scala 126:27]
  assign _GEN_3 = io_in_6_valid ? io_in_6_bits_idx : io_in_7_bits_idx; // @[Arbiter.scala 126:27]
  assign _GEN_4 = io_in_6_valid ? io_in_6_bits_addr : io_in_7_bits_addr; // @[Arbiter.scala 126:27]
  assign _GEN_13 = io_in_4_valid ? io_in_4_bits_data : _GEN_1; // @[Arbiter.scala 126:27]
  assign _GEN_14 = io_in_4_valid ? io_in_4_bits_way_en : _GEN_2; // @[Arbiter.scala 126:27]
  assign _GEN_15 = io_in_4_valid ? io_in_4_bits_idx : _GEN_3; // @[Arbiter.scala 126:27]
  assign _GEN_16 = io_in_4_valid ? io_in_4_bits_addr : _GEN_4; // @[Arbiter.scala 126:27]
  assign _GEN_19 = io_in_3_valid ? io_in_3_bits_data : _GEN_13; // @[Arbiter.scala 126:27]
  assign _GEN_20 = io_in_3_valid ? io_in_3_bits_way_en : _GEN_14; // @[Arbiter.scala 126:27]
  assign _GEN_21 = io_in_3_valid ? io_in_3_bits_idx : _GEN_15; // @[Arbiter.scala 126:27]
  assign _GEN_22 = io_in_3_valid ? io_in_3_bits_addr : _GEN_16; // @[Arbiter.scala 126:27]
  assign _GEN_23 = io_in_3_valid | io_in_4_valid; // @[Arbiter.scala 126:27]
  assign _GEN_25 = io_in_2_valid ? io_in_2_bits_data : _GEN_19; // @[Arbiter.scala 126:27]
  assign _GEN_26 = io_in_2_valid ? io_in_2_bits_way_en : _GEN_20; // @[Arbiter.scala 126:27]
  assign _GEN_27 = io_in_2_valid ? io_in_2_bits_idx : _GEN_21; // @[Arbiter.scala 126:27]
  assign _GEN_28 = io_in_2_valid ? io_in_2_bits_addr : _GEN_22; // @[Arbiter.scala 126:27]
  assign _GEN_29 = io_in_2_valid | _GEN_23; // @[Arbiter.scala 126:27]
  assign _GEN_31 = io_in_1_valid ? io_in_1_bits_data : _GEN_25; // @[Arbiter.scala 126:27]
  assign _GEN_32 = io_in_1_valid ? 4'h0 : _GEN_26; // @[Arbiter.scala 126:27]
  assign _GEN_33 = io_in_1_valid ? io_in_1_bits_idx : _GEN_27; // @[Arbiter.scala 126:27]
  assign _GEN_34 = io_in_1_valid ? io_in_1_bits_addr : _GEN_28; // @[Arbiter.scala 126:27]
  assign _GEN_35 = io_in_1_valid | _GEN_29; // @[Arbiter.scala 126:27]
  assign _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  assign _T_1 = _T | io_in_2_valid; // @[Arbiter.scala 31:68]
  assign _T_2 = _T_1 | io_in_3_valid; // @[Arbiter.scala 31:68]
  assign _T_3 = _T_2 | io_in_4_valid; // @[Arbiter.scala 31:68]
  assign _T_5 = _T_3 | io_in_6_valid; // @[Arbiter.scala 31:68]
  assign grant_7 = ~_T_5; // @[Arbiter.scala 31:78]
  assign io_in_4_ready = ~_T_2; // @[Arbiter.scala 134:14]
  assign io_in_5_ready = ~_T_3; // @[Arbiter.scala 134:14]
  assign io_in_6_ready = ~_T_3; // @[Arbiter.scala 134:14]
  assign io_in_7_ready = ~_T_5; // @[Arbiter.scala 134:14]
  assign io_out_valid = ~grant_7 | io_in_7_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_write = io_in_0_valid | _GEN_35; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_34; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_idx = io_in_0_valid ? io_in_0_bits_idx : _GEN_33; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_way_en = io_in_0_valid ? 4'hf : _GEN_32; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : _GEN_31; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign DCacheModuleImpl_Anon_1_covSum = 30'h0;
  assign io_covSum = DCacheModuleImpl_Anon_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module DCacheDataArray(
  input         clock,
  input         io_req_valid,
  input  [11:0] io_req_bits_addr,
  input         io_req_bits_write,
  input  [63:0] io_req_bits_wdata,
  input  [7:0]  io_req_bits_eccMask,
  input  [3:0]  io_req_bits_way_en,
  output [63:0] io_resp_0,
  output [63:0] io_resp_1,
  output [63:0] io_resp_2,
  output [63:0] io_resp_3,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [7:0] data_arrays_0_0 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_0;
  wire [7:0] data_arrays_0_0__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_0__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_0__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_0__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_0__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_0__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_0__T_51_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [8:0] data_arrays_0_0__T_51_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg [7:0] data_arrays_0_1 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_3;
  wire [7:0] data_arrays_0_1__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_1__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_1__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_1__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_1__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_1__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_1__T_51_en_pipe_0;
  reg [31:0] _RAND_4;
  reg [8:0] data_arrays_0_1__T_51_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [7:0] data_arrays_0_2 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_6;
  wire [7:0] data_arrays_0_2__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_2__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_2__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_2__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_2__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_2__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_2__T_51_en_pipe_0;
  reg [31:0] _RAND_7;
  reg [8:0] data_arrays_0_2__T_51_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [7:0] data_arrays_0_3 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_9;
  wire [7:0] data_arrays_0_3__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_3__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_3__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_3__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_3__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_3__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_3__T_51_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [8:0] data_arrays_0_3__T_51_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [7:0] data_arrays_0_4 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_12;
  wire [7:0] data_arrays_0_4__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_4__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_4__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_4__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_4__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_4__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_4__T_51_en_pipe_0;
  reg [31:0] _RAND_13;
  reg [8:0] data_arrays_0_4__T_51_addr_pipe_0;
  reg [31:0] _RAND_14;
  reg [7:0] data_arrays_0_5 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_15;
  wire [7:0] data_arrays_0_5__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_5__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_5__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_5__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_5__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_5__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_5__T_51_en_pipe_0;
  reg [31:0] _RAND_16;
  reg [8:0] data_arrays_0_5__T_51_addr_pipe_0;
  reg [31:0] _RAND_17;
  reg [7:0] data_arrays_0_6 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_18;
  wire [7:0] data_arrays_0_6__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_6__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_6__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_6__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_6__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_6__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_6__T_51_en_pipe_0;
  reg [31:0] _RAND_19;
  reg [8:0] data_arrays_0_6__T_51_addr_pipe_0;
  reg [31:0] _RAND_20;
  reg [7:0] data_arrays_0_7 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_21;
  wire [7:0] data_arrays_0_7__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_7__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_7__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_7__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_7__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_7__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_7__T_51_en_pipe_0;
  reg [31:0] _RAND_22;
  reg [8:0] data_arrays_0_7__T_51_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [7:0] data_arrays_0_8 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_24;
  wire [7:0] data_arrays_0_8__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_8__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_8__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_8__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_8__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_8__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_8__T_51_en_pipe_0;
  reg [31:0] _RAND_25;
  reg [8:0] data_arrays_0_8__T_51_addr_pipe_0;
  reg [31:0] _RAND_26;
  reg [7:0] data_arrays_0_9 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_27;
  wire [7:0] data_arrays_0_9__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_9__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_9__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_9__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_9__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_9__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_9__T_51_en_pipe_0;
  reg [31:0] _RAND_28;
  reg [8:0] data_arrays_0_9__T_51_addr_pipe_0;
  reg [31:0] _RAND_29;
  reg [7:0] data_arrays_0_10 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_30;
  wire [7:0] data_arrays_0_10__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_10__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_10__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_10__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_10__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_10__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_10__T_51_en_pipe_0;
  reg [31:0] _RAND_31;
  reg [8:0] data_arrays_0_10__T_51_addr_pipe_0;
  reg [31:0] _RAND_32;
  reg [7:0] data_arrays_0_11 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_33;
  wire [7:0] data_arrays_0_11__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_11__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_11__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_11__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_11__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_11__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_11__T_51_en_pipe_0;
  reg [31:0] _RAND_34;
  reg [8:0] data_arrays_0_11__T_51_addr_pipe_0;
  reg [31:0] _RAND_35;
  reg [7:0] data_arrays_0_12 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_36;
  wire [7:0] data_arrays_0_12__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_12__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_12__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_12__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_12__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_12__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_12__T_51_en_pipe_0;
  reg [31:0] _RAND_37;
  reg [8:0] data_arrays_0_12__T_51_addr_pipe_0;
  reg [31:0] _RAND_38;
  reg [7:0] data_arrays_0_13 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_39;
  wire [7:0] data_arrays_0_13__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_13__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_13__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_13__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_13__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_13__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_13__T_51_en_pipe_0;
  reg [31:0] _RAND_40;
  reg [8:0] data_arrays_0_13__T_51_addr_pipe_0;
  reg [31:0] _RAND_41;
  reg [7:0] data_arrays_0_14 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_42;
  wire [7:0] data_arrays_0_14__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_14__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_14__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_14__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_14__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_14__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_14__T_51_en_pipe_0;
  reg [31:0] _RAND_43;
  reg [8:0] data_arrays_0_14__T_51_addr_pipe_0;
  reg [31:0] _RAND_44;
  reg [7:0] data_arrays_0_15 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_45;
  wire [7:0] data_arrays_0_15__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_15__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_15__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_15__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_15__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_15__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_15__T_51_en_pipe_0;
  reg [31:0] _RAND_46;
  reg [8:0] data_arrays_0_15__T_51_addr_pipe_0;
  reg [31:0] _RAND_47;
  reg [7:0] data_arrays_0_16 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_48;
  wire [7:0] data_arrays_0_16__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_16__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_16__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_16__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_16__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_16__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_16__T_51_en_pipe_0;
  reg [31:0] _RAND_49;
  reg [8:0] data_arrays_0_16__T_51_addr_pipe_0;
  reg [31:0] _RAND_50;
  reg [7:0] data_arrays_0_17 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_51;
  wire [7:0] data_arrays_0_17__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_17__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_17__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_17__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_17__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_17__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_17__T_51_en_pipe_0;
  reg [31:0] _RAND_52;
  reg [8:0] data_arrays_0_17__T_51_addr_pipe_0;
  reg [31:0] _RAND_53;
  reg [7:0] data_arrays_0_18 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_54;
  wire [7:0] data_arrays_0_18__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_18__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_18__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_18__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_18__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_18__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_18__T_51_en_pipe_0;
  reg [31:0] _RAND_55;
  reg [8:0] data_arrays_0_18__T_51_addr_pipe_0;
  reg [31:0] _RAND_56;
  reg [7:0] data_arrays_0_19 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_57;
  wire [7:0] data_arrays_0_19__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_19__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_19__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_19__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_19__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_19__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_19__T_51_en_pipe_0;
  reg [31:0] _RAND_58;
  reg [8:0] data_arrays_0_19__T_51_addr_pipe_0;
  reg [31:0] _RAND_59;
  reg [7:0] data_arrays_0_20 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_60;
  wire [7:0] data_arrays_0_20__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_20__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_20__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_20__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_20__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_20__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_20__T_51_en_pipe_0;
  reg [31:0] _RAND_61;
  reg [8:0] data_arrays_0_20__T_51_addr_pipe_0;
  reg [31:0] _RAND_62;
  reg [7:0] data_arrays_0_21 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_63;
  wire [7:0] data_arrays_0_21__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_21__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_21__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_21__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_21__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_21__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_21__T_51_en_pipe_0;
  reg [31:0] _RAND_64;
  reg [8:0] data_arrays_0_21__T_51_addr_pipe_0;
  reg [31:0] _RAND_65;
  reg [7:0] data_arrays_0_22 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_66;
  wire [7:0] data_arrays_0_22__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_22__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_22__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_22__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_22__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_22__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_22__T_51_en_pipe_0;
  reg [31:0] _RAND_67;
  reg [8:0] data_arrays_0_22__T_51_addr_pipe_0;
  reg [31:0] _RAND_68;
  reg [7:0] data_arrays_0_23 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_69;
  wire [7:0] data_arrays_0_23__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_23__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_23__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_23__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_23__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_23__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_23__T_51_en_pipe_0;
  reg [31:0] _RAND_70;
  reg [8:0] data_arrays_0_23__T_51_addr_pipe_0;
  reg [31:0] _RAND_71;
  reg [7:0] data_arrays_0_24 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_72;
  wire [7:0] data_arrays_0_24__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_24__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_24__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_24__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_24__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_24__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_24__T_51_en_pipe_0;
  reg [31:0] _RAND_73;
  reg [8:0] data_arrays_0_24__T_51_addr_pipe_0;
  reg [31:0] _RAND_74;
  reg [7:0] data_arrays_0_25 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_75;
  wire [7:0] data_arrays_0_25__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_25__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_25__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_25__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_25__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_25__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_25__T_51_en_pipe_0;
  reg [31:0] _RAND_76;
  reg [8:0] data_arrays_0_25__T_51_addr_pipe_0;
  reg [31:0] _RAND_77;
  reg [7:0] data_arrays_0_26 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_78;
  wire [7:0] data_arrays_0_26__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_26__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_26__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_26__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_26__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_26__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_26__T_51_en_pipe_0;
  reg [31:0] _RAND_79;
  reg [8:0] data_arrays_0_26__T_51_addr_pipe_0;
  reg [31:0] _RAND_80;
  reg [7:0] data_arrays_0_27 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_81;
  wire [7:0] data_arrays_0_27__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_27__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_27__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_27__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_27__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_27__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_27__T_51_en_pipe_0;
  reg [31:0] _RAND_82;
  reg [8:0] data_arrays_0_27__T_51_addr_pipe_0;
  reg [31:0] _RAND_83;
  reg [7:0] data_arrays_0_28 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_84;
  wire [7:0] data_arrays_0_28__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_28__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_28__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_28__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_28__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_28__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_28__T_51_en_pipe_0;
  reg [31:0] _RAND_85;
  reg [8:0] data_arrays_0_28__T_51_addr_pipe_0;
  reg [31:0] _RAND_86;
  reg [7:0] data_arrays_0_29 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_87;
  wire [7:0] data_arrays_0_29__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_29__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_29__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_29__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_29__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_29__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_29__T_51_en_pipe_0;
  reg [31:0] _RAND_88;
  reg [8:0] data_arrays_0_29__T_51_addr_pipe_0;
  reg [31:0] _RAND_89;
  reg [7:0] data_arrays_0_30 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_90;
  wire [7:0] data_arrays_0_30__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_30__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_30__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_30__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_30__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_30__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_30__T_51_en_pipe_0;
  reg [31:0] _RAND_91;
  reg [8:0] data_arrays_0_30__T_51_addr_pipe_0;
  reg [31:0] _RAND_92;
  reg [7:0] data_arrays_0_31 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_93;
  wire [7:0] data_arrays_0_31__T_51_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_31__T_51_addr; // @[DescribedSRAM.scala 23:26]
  wire [7:0] data_arrays_0_31__T_45_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_31__T_45_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_31__T_45_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_31__T_45_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_31__T_51_en_pipe_0;
  reg [31:0] _RAND_94;
  reg [8:0] data_arrays_0_31__T_51_addr_pipe_0;
  reg [31:0] _RAND_95;
  wire  eccMask_0; // @[DCache.scala 50:79]
  wire  eccMask_1; // @[DCache.scala 50:79]
  wire  eccMask_2; // @[DCache.scala 50:79]
  wire  eccMask_3; // @[DCache.scala 50:79]
  wire  eccMask_4; // @[DCache.scala 50:79]
  wire  eccMask_5; // @[DCache.scala 50:79]
  wire  eccMask_6; // @[DCache.scala 50:79]
  wire  eccMask_7; // @[DCache.scala 50:79]
  wire [31:0] _T_54; // @[Cat.scala 29:58]
  wire [31:0] _T_57; // @[Cat.scala 29:58]
  wire [31:0] _T_60; // @[Cat.scala 29:58]
  wire [31:0] _T_63; // @[Cat.scala 29:58]
  wire [31:0] _T_66; // @[Cat.scala 29:58]
  wire [31:0] _T_69; // @[Cat.scala 29:58]
  wire [31:0] _T_72; // @[Cat.scala 29:58]
  wire [31:0] _T_75; // @[Cat.scala 29:58]
  wire [29:0] DCacheDataArray_covSum;
  assign data_arrays_0_0__T_51_addr = data_arrays_0_0__T_51_addr_pipe_0;
  assign data_arrays_0_0__T_51_data = data_arrays_0_0[data_arrays_0_0__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_0__T_45_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_0__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_0__T_45_mask = eccMask_0 & io_req_bits_way_en[0];
  assign data_arrays_0_0__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_1__T_51_addr = data_arrays_0_1__T_51_addr_pipe_0;
  assign data_arrays_0_1__T_51_data = data_arrays_0_1[data_arrays_0_1__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_1__T_45_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_1__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_1__T_45_mask = eccMask_1 & io_req_bits_way_en[0];
  assign data_arrays_0_1__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_2__T_51_addr = data_arrays_0_2__T_51_addr_pipe_0;
  assign data_arrays_0_2__T_51_data = data_arrays_0_2[data_arrays_0_2__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_2__T_45_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_2__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_2__T_45_mask = eccMask_2 & io_req_bits_way_en[0];
  assign data_arrays_0_2__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_3__T_51_addr = data_arrays_0_3__T_51_addr_pipe_0;
  assign data_arrays_0_3__T_51_data = data_arrays_0_3[data_arrays_0_3__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_3__T_45_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_3__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_3__T_45_mask = eccMask_3 & io_req_bits_way_en[0];
  assign data_arrays_0_3__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_4__T_51_addr = data_arrays_0_4__T_51_addr_pipe_0;
  assign data_arrays_0_4__T_51_data = data_arrays_0_4[data_arrays_0_4__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_4__T_45_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_4__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_4__T_45_mask = eccMask_4 & io_req_bits_way_en[0];
  assign data_arrays_0_4__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_5__T_51_addr = data_arrays_0_5__T_51_addr_pipe_0;
  assign data_arrays_0_5__T_51_data = data_arrays_0_5[data_arrays_0_5__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_5__T_45_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_5__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_5__T_45_mask = eccMask_5 & io_req_bits_way_en[0];
  assign data_arrays_0_5__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_6__T_51_addr = data_arrays_0_6__T_51_addr_pipe_0;
  assign data_arrays_0_6__T_51_data = data_arrays_0_6[data_arrays_0_6__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_6__T_45_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_6__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_6__T_45_mask = eccMask_6 & io_req_bits_way_en[0];
  assign data_arrays_0_6__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_7__T_51_addr = data_arrays_0_7__T_51_addr_pipe_0;
  assign data_arrays_0_7__T_51_data = data_arrays_0_7[data_arrays_0_7__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_7__T_45_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_7__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_7__T_45_mask = eccMask_7 & io_req_bits_way_en[0];
  assign data_arrays_0_7__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_8__T_51_addr = data_arrays_0_8__T_51_addr_pipe_0;
  assign data_arrays_0_8__T_51_data = data_arrays_0_8[data_arrays_0_8__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_8__T_45_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_8__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_8__T_45_mask = eccMask_0 & io_req_bits_way_en[1];
  assign data_arrays_0_8__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_9__T_51_addr = data_arrays_0_9__T_51_addr_pipe_0;
  assign data_arrays_0_9__T_51_data = data_arrays_0_9[data_arrays_0_9__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_9__T_45_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_9__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_9__T_45_mask = eccMask_1 & io_req_bits_way_en[1];
  assign data_arrays_0_9__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_10__T_51_addr = data_arrays_0_10__T_51_addr_pipe_0;
  assign data_arrays_0_10__T_51_data = data_arrays_0_10[data_arrays_0_10__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_10__T_45_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_10__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_10__T_45_mask = eccMask_2 & io_req_bits_way_en[1];
  assign data_arrays_0_10__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_11__T_51_addr = data_arrays_0_11__T_51_addr_pipe_0;
  assign data_arrays_0_11__T_51_data = data_arrays_0_11[data_arrays_0_11__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_11__T_45_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_11__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_11__T_45_mask = eccMask_3 & io_req_bits_way_en[1];
  assign data_arrays_0_11__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_12__T_51_addr = data_arrays_0_12__T_51_addr_pipe_0;
  assign data_arrays_0_12__T_51_data = data_arrays_0_12[data_arrays_0_12__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_12__T_45_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_12__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_12__T_45_mask = eccMask_4 & io_req_bits_way_en[1];
  assign data_arrays_0_12__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_13__T_51_addr = data_arrays_0_13__T_51_addr_pipe_0;
  assign data_arrays_0_13__T_51_data = data_arrays_0_13[data_arrays_0_13__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_13__T_45_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_13__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_13__T_45_mask = eccMask_5 & io_req_bits_way_en[1];
  assign data_arrays_0_13__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_14__T_51_addr = data_arrays_0_14__T_51_addr_pipe_0;
  assign data_arrays_0_14__T_51_data = data_arrays_0_14[data_arrays_0_14__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_14__T_45_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_14__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_14__T_45_mask = eccMask_6 & io_req_bits_way_en[1];
  assign data_arrays_0_14__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_15__T_51_addr = data_arrays_0_15__T_51_addr_pipe_0;
  assign data_arrays_0_15__T_51_data = data_arrays_0_15[data_arrays_0_15__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_15__T_45_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_15__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_15__T_45_mask = eccMask_7 & io_req_bits_way_en[1];
  assign data_arrays_0_15__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_16__T_51_addr = data_arrays_0_16__T_51_addr_pipe_0;
  assign data_arrays_0_16__T_51_data = data_arrays_0_16[data_arrays_0_16__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_16__T_45_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_16__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_16__T_45_mask = eccMask_0 & io_req_bits_way_en[2];
  assign data_arrays_0_16__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_17__T_51_addr = data_arrays_0_17__T_51_addr_pipe_0;
  assign data_arrays_0_17__T_51_data = data_arrays_0_17[data_arrays_0_17__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_17__T_45_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_17__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_17__T_45_mask = eccMask_1 & io_req_bits_way_en[2];
  assign data_arrays_0_17__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_18__T_51_addr = data_arrays_0_18__T_51_addr_pipe_0;
  assign data_arrays_0_18__T_51_data = data_arrays_0_18[data_arrays_0_18__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_18__T_45_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_18__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_18__T_45_mask = eccMask_2 & io_req_bits_way_en[2];
  assign data_arrays_0_18__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_19__T_51_addr = data_arrays_0_19__T_51_addr_pipe_0;
  assign data_arrays_0_19__T_51_data = data_arrays_0_19[data_arrays_0_19__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_19__T_45_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_19__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_19__T_45_mask = eccMask_3 & io_req_bits_way_en[2];
  assign data_arrays_0_19__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_20__T_51_addr = data_arrays_0_20__T_51_addr_pipe_0;
  assign data_arrays_0_20__T_51_data = data_arrays_0_20[data_arrays_0_20__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_20__T_45_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_20__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_20__T_45_mask = eccMask_4 & io_req_bits_way_en[2];
  assign data_arrays_0_20__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_21__T_51_addr = data_arrays_0_21__T_51_addr_pipe_0;
  assign data_arrays_0_21__T_51_data = data_arrays_0_21[data_arrays_0_21__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_21__T_45_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_21__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_21__T_45_mask = eccMask_5 & io_req_bits_way_en[2];
  assign data_arrays_0_21__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_22__T_51_addr = data_arrays_0_22__T_51_addr_pipe_0;
  assign data_arrays_0_22__T_51_data = data_arrays_0_22[data_arrays_0_22__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_22__T_45_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_22__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_22__T_45_mask = eccMask_6 & io_req_bits_way_en[2];
  assign data_arrays_0_22__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_23__T_51_addr = data_arrays_0_23__T_51_addr_pipe_0;
  assign data_arrays_0_23__T_51_data = data_arrays_0_23[data_arrays_0_23__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_23__T_45_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_23__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_23__T_45_mask = eccMask_7 & io_req_bits_way_en[2];
  assign data_arrays_0_23__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_24__T_51_addr = data_arrays_0_24__T_51_addr_pipe_0;
  assign data_arrays_0_24__T_51_data = data_arrays_0_24[data_arrays_0_24__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_24__T_45_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_24__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_24__T_45_mask = eccMask_0 & io_req_bits_way_en[3];
  assign data_arrays_0_24__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_25__T_51_addr = data_arrays_0_25__T_51_addr_pipe_0;
  assign data_arrays_0_25__T_51_data = data_arrays_0_25[data_arrays_0_25__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_25__T_45_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_25__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_25__T_45_mask = eccMask_1 & io_req_bits_way_en[3];
  assign data_arrays_0_25__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_26__T_51_addr = data_arrays_0_26__T_51_addr_pipe_0;
  assign data_arrays_0_26__T_51_data = data_arrays_0_26[data_arrays_0_26__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_26__T_45_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_26__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_26__T_45_mask = eccMask_2 & io_req_bits_way_en[3];
  assign data_arrays_0_26__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_27__T_51_addr = data_arrays_0_27__T_51_addr_pipe_0;
  assign data_arrays_0_27__T_51_data = data_arrays_0_27[data_arrays_0_27__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_27__T_45_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_27__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_27__T_45_mask = eccMask_3 & io_req_bits_way_en[3];
  assign data_arrays_0_27__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_28__T_51_addr = data_arrays_0_28__T_51_addr_pipe_0;
  assign data_arrays_0_28__T_51_data = data_arrays_0_28[data_arrays_0_28__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_28__T_45_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_28__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_28__T_45_mask = eccMask_4 & io_req_bits_way_en[3];
  assign data_arrays_0_28__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_29__T_51_addr = data_arrays_0_29__T_51_addr_pipe_0;
  assign data_arrays_0_29__T_51_data = data_arrays_0_29[data_arrays_0_29__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_29__T_45_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_29__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_29__T_45_mask = eccMask_5 & io_req_bits_way_en[3];
  assign data_arrays_0_29__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_30__T_51_addr = data_arrays_0_30__T_51_addr_pipe_0;
  assign data_arrays_0_30__T_51_data = data_arrays_0_30[data_arrays_0_30__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_30__T_45_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_30__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_30__T_45_mask = eccMask_6 & io_req_bits_way_en[3];
  assign data_arrays_0_30__T_45_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_31__T_51_addr = data_arrays_0_31__T_51_addr_pipe_0;
  assign data_arrays_0_31__T_51_data = data_arrays_0_31[data_arrays_0_31__T_51_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_31__T_45_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_31__T_45_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_31__T_45_mask = eccMask_7 & io_req_bits_way_en[3];
  assign data_arrays_0_31__T_45_en = io_req_valid & io_req_bits_write;
  assign eccMask_0 = io_req_bits_eccMask[0]; // @[DCache.scala 50:79]
  assign eccMask_1 = io_req_bits_eccMask[1]; // @[DCache.scala 50:79]
  assign eccMask_2 = io_req_bits_eccMask[2]; // @[DCache.scala 50:79]
  assign eccMask_3 = io_req_bits_eccMask[3]; // @[DCache.scala 50:79]
  assign eccMask_4 = io_req_bits_eccMask[4]; // @[DCache.scala 50:79]
  assign eccMask_5 = io_req_bits_eccMask[5]; // @[DCache.scala 50:79]
  assign eccMask_6 = io_req_bits_eccMask[6]; // @[DCache.scala 50:79]
  assign eccMask_7 = io_req_bits_eccMask[7]; // @[DCache.scala 50:79]
  assign _T_54 = {data_arrays_0_3__T_51_data,data_arrays_0_2__T_51_data,data_arrays_0_1__T_51_data,data_arrays_0_0__T_51_data}; // @[Cat.scala 29:58]
  assign _T_57 = {data_arrays_0_7__T_51_data,data_arrays_0_6__T_51_data,data_arrays_0_5__T_51_data,data_arrays_0_4__T_51_data}; // @[Cat.scala 29:58]
  assign _T_60 = {data_arrays_0_11__T_51_data,data_arrays_0_10__T_51_data,data_arrays_0_9__T_51_data,data_arrays_0_8__T_51_data}; // @[Cat.scala 29:58]
  assign _T_63 = {data_arrays_0_15__T_51_data,data_arrays_0_14__T_51_data,data_arrays_0_13__T_51_data,data_arrays_0_12__T_51_data}; // @[Cat.scala 29:58]
  assign _T_66 = {data_arrays_0_19__T_51_data,data_arrays_0_18__T_51_data,data_arrays_0_17__T_51_data,data_arrays_0_16__T_51_data}; // @[Cat.scala 29:58]
  assign _T_69 = {data_arrays_0_23__T_51_data,data_arrays_0_22__T_51_data,data_arrays_0_21__T_51_data,data_arrays_0_20__T_51_data}; // @[Cat.scala 29:58]
  assign _T_72 = {data_arrays_0_27__T_51_data,data_arrays_0_26__T_51_data,data_arrays_0_25__T_51_data,data_arrays_0_24__T_51_data}; // @[Cat.scala 29:58]
  assign _T_75 = {data_arrays_0_31__T_51_data,data_arrays_0_30__T_51_data,data_arrays_0_29__T_51_data,data_arrays_0_28__T_51_data}; // @[Cat.scala 29:58]
  assign io_resp_0 = {_T_57,_T_54}; // @[DCache.scala 73:69]
  assign io_resp_1 = {_T_63,_T_60}; // @[DCache.scala 73:69]
  assign io_resp_2 = {_T_69,_T_66}; // @[DCache.scala 73:69]
  assign io_resp_3 = {_T_75,_T_72}; // @[DCache.scala 73:69]
  assign DCacheDataArray_covSum = 30'h0;
  assign io_covSum = DCacheDataArray_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_0[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  data_arrays_0_0__T_51_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  data_arrays_0_0__T_51_addr_pipe_0 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_1[initvar] = _RAND_3[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  data_arrays_0_1__T_51_en_pipe_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  data_arrays_0_1__T_51_addr_pipe_0 = _RAND_5[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_2[initvar] = _RAND_6[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_arrays_0_2__T_51_en_pipe_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  data_arrays_0_2__T_51_addr_pipe_0 = _RAND_8[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_3[initvar] = _RAND_9[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_arrays_0_3__T_51_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  data_arrays_0_3__T_51_addr_pipe_0 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_4[initvar] = _RAND_12[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  data_arrays_0_4__T_51_en_pipe_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  data_arrays_0_4__T_51_addr_pipe_0 = _RAND_14[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_5[initvar] = _RAND_15[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  data_arrays_0_5__T_51_en_pipe_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  data_arrays_0_5__T_51_addr_pipe_0 = _RAND_17[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_6[initvar] = _RAND_18[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  data_arrays_0_6__T_51_en_pipe_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  data_arrays_0_6__T_51_addr_pipe_0 = _RAND_20[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_7[initvar] = _RAND_21[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  data_arrays_0_7__T_51_en_pipe_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  data_arrays_0_7__T_51_addr_pipe_0 = _RAND_23[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_8[initvar] = _RAND_24[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  data_arrays_0_8__T_51_en_pipe_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  data_arrays_0_8__T_51_addr_pipe_0 = _RAND_26[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_9[initvar] = _RAND_27[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  data_arrays_0_9__T_51_en_pipe_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  data_arrays_0_9__T_51_addr_pipe_0 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_10[initvar] = _RAND_30[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  data_arrays_0_10__T_51_en_pipe_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  data_arrays_0_10__T_51_addr_pipe_0 = _RAND_32[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_11[initvar] = _RAND_33[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  data_arrays_0_11__T_51_en_pipe_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  data_arrays_0_11__T_51_addr_pipe_0 = _RAND_35[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_12[initvar] = _RAND_36[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  data_arrays_0_12__T_51_en_pipe_0 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  data_arrays_0_12__T_51_addr_pipe_0 = _RAND_38[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_13[initvar] = _RAND_39[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  data_arrays_0_13__T_51_en_pipe_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  data_arrays_0_13__T_51_addr_pipe_0 = _RAND_41[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_14[initvar] = _RAND_42[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  data_arrays_0_14__T_51_en_pipe_0 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  data_arrays_0_14__T_51_addr_pipe_0 = _RAND_44[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_15[initvar] = _RAND_45[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  data_arrays_0_15__T_51_en_pipe_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  data_arrays_0_15__T_51_addr_pipe_0 = _RAND_47[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_16[initvar] = _RAND_48[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  data_arrays_0_16__T_51_en_pipe_0 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  data_arrays_0_16__T_51_addr_pipe_0 = _RAND_50[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_17[initvar] = _RAND_51[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  data_arrays_0_17__T_51_en_pipe_0 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  data_arrays_0_17__T_51_addr_pipe_0 = _RAND_53[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_18[initvar] = _RAND_54[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  data_arrays_0_18__T_51_en_pipe_0 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  data_arrays_0_18__T_51_addr_pipe_0 = _RAND_56[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_19[initvar] = _RAND_57[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  data_arrays_0_19__T_51_en_pipe_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  data_arrays_0_19__T_51_addr_pipe_0 = _RAND_59[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_20[initvar] = _RAND_60[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  data_arrays_0_20__T_51_en_pipe_0 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  data_arrays_0_20__T_51_addr_pipe_0 = _RAND_62[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_21[initvar] = _RAND_63[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  data_arrays_0_21__T_51_en_pipe_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  data_arrays_0_21__T_51_addr_pipe_0 = _RAND_65[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_22[initvar] = _RAND_66[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  data_arrays_0_22__T_51_en_pipe_0 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  data_arrays_0_22__T_51_addr_pipe_0 = _RAND_68[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_23[initvar] = _RAND_69[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  data_arrays_0_23__T_51_en_pipe_0 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  data_arrays_0_23__T_51_addr_pipe_0 = _RAND_71[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_24[initvar] = _RAND_72[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  data_arrays_0_24__T_51_en_pipe_0 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  data_arrays_0_24__T_51_addr_pipe_0 = _RAND_74[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_25[initvar] = _RAND_75[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  data_arrays_0_25__T_51_en_pipe_0 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  data_arrays_0_25__T_51_addr_pipe_0 = _RAND_77[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_26[initvar] = _RAND_78[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  data_arrays_0_26__T_51_en_pipe_0 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  data_arrays_0_26__T_51_addr_pipe_0 = _RAND_80[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_27[initvar] = _RAND_81[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  data_arrays_0_27__T_51_en_pipe_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  data_arrays_0_27__T_51_addr_pipe_0 = _RAND_83[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_28[initvar] = _RAND_84[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  data_arrays_0_28__T_51_en_pipe_0 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  data_arrays_0_28__T_51_addr_pipe_0 = _RAND_86[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_29[initvar] = _RAND_87[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  data_arrays_0_29__T_51_en_pipe_0 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  data_arrays_0_29__T_51_addr_pipe_0 = _RAND_89[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_30[initvar] = _RAND_90[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  data_arrays_0_30__T_51_en_pipe_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  data_arrays_0_30__T_51_addr_pipe_0 = _RAND_92[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_31[initvar] = _RAND_93[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  data_arrays_0_31__T_51_en_pipe_0 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  data_arrays_0_31__T_51_addr_pipe_0 = _RAND_95[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(data_arrays_0_0__T_45_en & data_arrays_0_0__T_45_mask) begin
      data_arrays_0_0[data_arrays_0_0__T_45_addr] <= data_arrays_0_0__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_0__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_0__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_0__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_0__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_1__T_45_en & data_arrays_0_1__T_45_mask) begin
      data_arrays_0_1[data_arrays_0_1__T_45_addr] <= data_arrays_0_1__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_1__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_1__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_1__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_1__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_2__T_45_en & data_arrays_0_2__T_45_mask) begin
      data_arrays_0_2[data_arrays_0_2__T_45_addr] <= data_arrays_0_2__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_2__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_2__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_2__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_2__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_3__T_45_en & data_arrays_0_3__T_45_mask) begin
      data_arrays_0_3[data_arrays_0_3__T_45_addr] <= data_arrays_0_3__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_3__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_3__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_3__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_3__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_4__T_45_en & data_arrays_0_4__T_45_mask) begin
      data_arrays_0_4[data_arrays_0_4__T_45_addr] <= data_arrays_0_4__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_4__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_4__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_4__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_4__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_5__T_45_en & data_arrays_0_5__T_45_mask) begin
      data_arrays_0_5[data_arrays_0_5__T_45_addr] <= data_arrays_0_5__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_5__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_5__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_5__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_5__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_6__T_45_en & data_arrays_0_6__T_45_mask) begin
      data_arrays_0_6[data_arrays_0_6__T_45_addr] <= data_arrays_0_6__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_6__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_6__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_6__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_6__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_7__T_45_en & data_arrays_0_7__T_45_mask) begin
      data_arrays_0_7[data_arrays_0_7__T_45_addr] <= data_arrays_0_7__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_7__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_7__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_7__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_7__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_8__T_45_en & data_arrays_0_8__T_45_mask) begin
      data_arrays_0_8[data_arrays_0_8__T_45_addr] <= data_arrays_0_8__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_8__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_8__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_8__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_8__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_9__T_45_en & data_arrays_0_9__T_45_mask) begin
      data_arrays_0_9[data_arrays_0_9__T_45_addr] <= data_arrays_0_9__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_9__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_9__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_9__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_9__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_10__T_45_en & data_arrays_0_10__T_45_mask) begin
      data_arrays_0_10[data_arrays_0_10__T_45_addr] <= data_arrays_0_10__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_10__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_10__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_10__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_10__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_11__T_45_en & data_arrays_0_11__T_45_mask) begin
      data_arrays_0_11[data_arrays_0_11__T_45_addr] <= data_arrays_0_11__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_11__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_11__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_11__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_11__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_12__T_45_en & data_arrays_0_12__T_45_mask) begin
      data_arrays_0_12[data_arrays_0_12__T_45_addr] <= data_arrays_0_12__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_12__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_12__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_12__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_12__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_13__T_45_en & data_arrays_0_13__T_45_mask) begin
      data_arrays_0_13[data_arrays_0_13__T_45_addr] <= data_arrays_0_13__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_13__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_13__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_13__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_13__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_14__T_45_en & data_arrays_0_14__T_45_mask) begin
      data_arrays_0_14[data_arrays_0_14__T_45_addr] <= data_arrays_0_14__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_14__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_14__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_14__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_14__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_15__T_45_en & data_arrays_0_15__T_45_mask) begin
      data_arrays_0_15[data_arrays_0_15__T_45_addr] <= data_arrays_0_15__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_15__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_15__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_15__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_15__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_16__T_45_en & data_arrays_0_16__T_45_mask) begin
      data_arrays_0_16[data_arrays_0_16__T_45_addr] <= data_arrays_0_16__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_16__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_16__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_16__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_16__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_17__T_45_en & data_arrays_0_17__T_45_mask) begin
      data_arrays_0_17[data_arrays_0_17__T_45_addr] <= data_arrays_0_17__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_17__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_17__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_17__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_17__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_18__T_45_en & data_arrays_0_18__T_45_mask) begin
      data_arrays_0_18[data_arrays_0_18__T_45_addr] <= data_arrays_0_18__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_18__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_18__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_18__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_18__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_19__T_45_en & data_arrays_0_19__T_45_mask) begin
      data_arrays_0_19[data_arrays_0_19__T_45_addr] <= data_arrays_0_19__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_19__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_19__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_19__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_19__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_20__T_45_en & data_arrays_0_20__T_45_mask) begin
      data_arrays_0_20[data_arrays_0_20__T_45_addr] <= data_arrays_0_20__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_20__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_20__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_20__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_20__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_21__T_45_en & data_arrays_0_21__T_45_mask) begin
      data_arrays_0_21[data_arrays_0_21__T_45_addr] <= data_arrays_0_21__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_21__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_21__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_21__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_21__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_22__T_45_en & data_arrays_0_22__T_45_mask) begin
      data_arrays_0_22[data_arrays_0_22__T_45_addr] <= data_arrays_0_22__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_22__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_22__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_22__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_22__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_23__T_45_en & data_arrays_0_23__T_45_mask) begin
      data_arrays_0_23[data_arrays_0_23__T_45_addr] <= data_arrays_0_23__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_23__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_23__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_23__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_23__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_24__T_45_en & data_arrays_0_24__T_45_mask) begin
      data_arrays_0_24[data_arrays_0_24__T_45_addr] <= data_arrays_0_24__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_24__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_24__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_24__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_24__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_25__T_45_en & data_arrays_0_25__T_45_mask) begin
      data_arrays_0_25[data_arrays_0_25__T_45_addr] <= data_arrays_0_25__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_25__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_25__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_25__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_25__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_26__T_45_en & data_arrays_0_26__T_45_mask) begin
      data_arrays_0_26[data_arrays_0_26__T_45_addr] <= data_arrays_0_26__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_26__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_26__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_26__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_26__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_27__T_45_en & data_arrays_0_27__T_45_mask) begin
      data_arrays_0_27[data_arrays_0_27__T_45_addr] <= data_arrays_0_27__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_27__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_27__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_27__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_27__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_28__T_45_en & data_arrays_0_28__T_45_mask) begin
      data_arrays_0_28[data_arrays_0_28__T_45_addr] <= data_arrays_0_28__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_28__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_28__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_28__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_28__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_29__T_45_en & data_arrays_0_29__T_45_mask) begin
      data_arrays_0_29[data_arrays_0_29__T_45_addr] <= data_arrays_0_29__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_29__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_29__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_29__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_29__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_30__T_45_en & data_arrays_0_30__T_45_mask) begin
      data_arrays_0_30[data_arrays_0_30__T_45_addr] <= data_arrays_0_30__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_30__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_30__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_30__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_30__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_31__T_45_en & data_arrays_0_31__T_45_mask) begin
      data_arrays_0_31[data_arrays_0_31__T_45_addr] <= data_arrays_0_31__T_45_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_31__T_51_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_31__T_51_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_31__T_51_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_31__T_51_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
  end
endmodule
module DCacheModuleImpl_Anon_2(
  input         io_in_0_valid,
  input  [11:0] io_in_0_bits_addr,
  input         io_in_0_bits_write,
  input  [63:0] io_in_0_bits_wdata,
  input  [7:0]  io_in_0_bits_eccMask,
  input  [3:0]  io_in_0_bits_way_en,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [11:0] io_in_1_bits_addr,
  input         io_in_1_bits_write,
  input  [63:0] io_in_1_bits_wdata,
  input  [7:0]  io_in_1_bits_eccMask,
  input  [3:0]  io_in_1_bits_way_en,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [11:0] io_in_2_bits_addr,
  input  [63:0] io_in_2_bits_wdata,
  input  [7:0]  io_in_2_bits_eccMask,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [11:0] io_in_3_bits_addr,
  input  [63:0] io_in_3_bits_wdata,
  input  [7:0]  io_in_3_bits_eccMask,
  output        io_out_valid,
  output [11:0] io_out_bits_addr,
  output        io_out_bits_write,
  output [63:0] io_out_bits_wdata,
  output [7:0]  io_out_bits_eccMask,
  output [3:0]  io_out_bits_way_en,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [7:0] _GEN_2; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_4; // @[Arbiter.scala 126:27]
  wire [11:0] _GEN_6; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_8; // @[Arbiter.scala 126:27]
  wire [7:0] _GEN_9; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_11; // @[Arbiter.scala 126:27]
  wire  _GEN_12; // @[Arbiter.scala 126:27]
  wire [11:0] _GEN_13; // @[Arbiter.scala 126:27]
  wire  _T; // @[Arbiter.scala 31:68]
  wire  _T_1; // @[Arbiter.scala 31:68]
  wire  grant_3; // @[Arbiter.scala 31:78]
  wire [29:0] DCacheModuleImpl_Anon_2_covSum;
  assign _GEN_2 = io_in_2_valid ? io_in_2_bits_eccMask : io_in_3_bits_eccMask; // @[Arbiter.scala 126:27]
  assign _GEN_4 = io_in_2_valid ? io_in_2_bits_wdata : io_in_3_bits_wdata; // @[Arbiter.scala 126:27]
  assign _GEN_6 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr; // @[Arbiter.scala 126:27]
  assign _GEN_8 = io_in_1_valid ? io_in_1_bits_way_en : 4'hf; // @[Arbiter.scala 126:27]
  assign _GEN_9 = io_in_1_valid ? 8'hff : _GEN_2; // @[Arbiter.scala 126:27]
  assign _GEN_11 = io_in_1_valid ? io_in_1_bits_wdata : _GEN_4; // @[Arbiter.scala 126:27]
  assign _GEN_12 = io_in_1_valid & io_in_1_bits_write; // @[Arbiter.scala 126:27]
  assign _GEN_13 = io_in_1_valid ? io_in_1_bits_addr : _GEN_6; // @[Arbiter.scala 126:27]
  assign _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  assign _T_1 = _T | io_in_2_valid; // @[Arbiter.scala 31:68]
  assign grant_3 = ~_T_1; // @[Arbiter.scala 31:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 134:14]
  assign io_in_2_ready = ~_T; // @[Arbiter.scala 134:14]
  assign io_in_3_ready = ~_T_1; // @[Arbiter.scala 134:14]
  assign io_out_valid = ~grant_3 | io_in_3_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_13; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_write = io_in_0_valid ? io_in_0_bits_write : _GEN_12; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : _GEN_11; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_eccMask = io_in_0_valid ? io_in_0_bits_eccMask : _GEN_9; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_way_en = io_in_0_valid ? io_in_0_bits_way_en : _GEN_8; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign DCacheModuleImpl_Anon_2_covSum = 30'h0;
  assign io_covSum = DCacheModuleImpl_Anon_2_covSum;
  assign metaAssert = 1'h0;
endmodule
module AMOALU(
  input  [7:0]  io_mask,
  input  [4:0]  io_cmd,
  input  [63:0] io_lhs,
  input  [63:0] io_rhs,
  output [63:0] io_out,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  _T; // @[AMOALU.scala 64:20]
  wire  _T_1; // @[AMOALU.scala 64:43]
  wire  max; // @[AMOALU.scala 64:33]
  wire  _T_2; // @[AMOALU.scala 65:20]
  wire  _T_3; // @[AMOALU.scala 65:43]
  wire  min; // @[AMOALU.scala 65:33]
  wire  add; // @[AMOALU.scala 66:20]
  wire  _T_4; // @[AMOALU.scala 67:26]
  wire  _T_5; // @[AMOALU.scala 67:48]
  wire  logic_and; // @[AMOALU.scala 67:38]
  wire  _T_6; // @[AMOALU.scala 68:26]
  wire  logic_xor; // @[AMOALU.scala 68:39]
  wire [31:0] _T_10; // @[AMOALU.scala 72:79]
  wire [63:0] _T_11; // @[AMOALU.scala 72:98]
  wire [63:0] _T_13; // @[AMOALU.scala 73:13]
  wire [63:0] _T_14; // @[AMOALU.scala 73:31]
  wire [63:0] adder_out; // @[AMOALU.scala 73:21]
  wire [4:0] _T_18; // @[AMOALU.scala 86:17]
  wire  _T_20; // @[AMOALU.scala 86:25]
  wire  _T_23; // @[AMOALU.scala 88:18]
  wire  _T_26; // @[AMOALU.scala 80:24]
  wire  _T_29; // @[AMOALU.scala 80:53]
  wire  _T_32; // @[AMOALU.scala 79:35]
  wire  _T_33; // @[AMOALU.scala 80:69]
  wire  _T_34; // @[AMOALU.scala 80:38]
  wire  _T_37; // @[AMOALU.scala 88:58]
  wire  _T_38; // @[AMOALU.scala 88:10]
  wire  _T_46; // @[AMOALU.scala 88:18]
  wire  _T_52; // @[AMOALU.scala 88:58]
  wire  _T_53; // @[AMOALU.scala 88:10]
  wire  less; // @[Mux.scala 47:69]
  wire  _T_54; // @[AMOALU.scala 94:23]
  wire [63:0] minmax; // @[AMOALU.scala 94:19]
  wire [63:0] _T_55; // @[AMOALU.scala 96:27]
  wire [63:0] _T_56; // @[AMOALU.scala 96:8]
  wire [63:0] _T_57; // @[AMOALU.scala 97:27]
  wire [63:0] _T_58; // @[AMOALU.scala 97:8]
  wire [63:0] logic_; // @[AMOALU.scala 96:42]
  wire  _T_59; // @[AMOALU.scala 100:19]
  wire [63:0] _T_60; // @[AMOALU.scala 100:8]
  wire [63:0] out; // @[AMOALU.scala 99:8]
  wire [7:0] _T_70; // @[Bitwise.scala 72:12]
  wire [7:0] _T_72; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76; // @[Bitwise.scala 72:12]
  wire [7:0] _T_78; // @[Bitwise.scala 72:12]
  wire [7:0] _T_80; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84; // @[Bitwise.scala 72:12]
  wire [63:0] wmask; // @[Cat.scala 29:58]
  wire [63:0] _T_91; // @[AMOALU.scala 104:19]
  wire [63:0] _T_93; // @[AMOALU.scala 104:34]
  wire [29:0] AMOALU_covSum;
  assign _T = io_cmd == 5'hd; // @[AMOALU.scala 64:20]
  assign _T_1 = io_cmd == 5'hf; // @[AMOALU.scala 64:43]
  assign max = _T | _T_1; // @[AMOALU.scala 64:33]
  assign _T_2 = io_cmd == 5'hc; // @[AMOALU.scala 65:20]
  assign _T_3 = io_cmd == 5'he; // @[AMOALU.scala 65:43]
  assign min = _T_2 | _T_3; // @[AMOALU.scala 65:33]
  assign add = io_cmd == 5'h8; // @[AMOALU.scala 66:20]
  assign _T_4 = io_cmd == 5'ha; // @[AMOALU.scala 67:26]
  assign _T_5 = io_cmd == 5'hb; // @[AMOALU.scala 67:48]
  assign logic_and = _T_4 | _T_5; // @[AMOALU.scala 67:38]
  assign _T_6 = io_cmd == 5'h9; // @[AMOALU.scala 68:26]
  assign logic_xor = _T_6 | _T_4; // @[AMOALU.scala 68:39]
  assign _T_10 = {~io_mask[3], 31'h0}; // @[AMOALU.scala 72:79]
  assign _T_11 = {{32'd0}, _T_10}; // @[AMOALU.scala 72:98]
  assign _T_13 = io_lhs & ~_T_11; // @[AMOALU.scala 73:13]
  assign _T_14 = io_rhs & ~_T_11; // @[AMOALU.scala 73:31]
  assign adder_out = _T_13 + _T_14; // @[AMOALU.scala 73:21]
  assign _T_18 = io_cmd & 5'h2; // @[AMOALU.scala 86:17]
  assign _T_20 = _T_18 == 5'h0; // @[AMOALU.scala 86:25]
  assign _T_23 = io_lhs[63] == io_rhs[63]; // @[AMOALU.scala 88:18]
  assign _T_26 = io_lhs[63:32] < io_rhs[63:32]; // @[AMOALU.scala 80:24]
  assign _T_29 = io_lhs[63:32] == io_rhs[63:32]; // @[AMOALU.scala 80:53]
  assign _T_32 = io_lhs[31:0] < io_rhs[31:0]; // @[AMOALU.scala 79:35]
  assign _T_33 = _T_29 & _T_32; // @[AMOALU.scala 80:69]
  assign _T_34 = _T_26 | _T_33; // @[AMOALU.scala 80:38]
  assign _T_37 = _T_20 ? io_lhs[63] : io_rhs[63]; // @[AMOALU.scala 88:58]
  assign _T_38 = _T_23 ? _T_34 : _T_37; // @[AMOALU.scala 88:10]
  assign _T_46 = io_lhs[31] == io_rhs[31]; // @[AMOALU.scala 88:18]
  assign _T_52 = _T_20 ? io_lhs[31] : io_rhs[31]; // @[AMOALU.scala 88:58]
  assign _T_53 = _T_46 ? _T_32 : _T_52; // @[AMOALU.scala 88:10]
  assign less = io_mask[4] ? _T_38 : _T_53; // @[Mux.scala 47:69]
  assign _T_54 = less ? min : max; // @[AMOALU.scala 94:23]
  assign minmax = _T_54 ? io_lhs : io_rhs; // @[AMOALU.scala 94:19]
  assign _T_55 = io_lhs & io_rhs; // @[AMOALU.scala 96:27]
  assign _T_56 = logic_and ? _T_55 : 64'h0; // @[AMOALU.scala 96:8]
  assign _T_57 = io_lhs ^ io_rhs; // @[AMOALU.scala 97:27]
  assign _T_58 = logic_xor ? _T_57 : 64'h0; // @[AMOALU.scala 97:8]
  assign logic_ = _T_56 | _T_58; // @[AMOALU.scala 96:42]
  assign _T_59 = logic_and | logic_xor; // @[AMOALU.scala 100:19]
  assign _T_60 = _T_59 ? logic_ : minmax; // @[AMOALU.scala 100:8]
  assign out = add ? adder_out : _T_60; // @[AMOALU.scala 99:8]
  assign _T_70 = io_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_72 = io_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_74 = io_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_76 = io_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_78 = io_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_80 = io_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_82 = io_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_84 = io_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign wmask = {_T_84,_T_82,_T_80,_T_78,_T_76,_T_74,_T_72,_T_70}; // @[Cat.scala 29:58]
  assign _T_91 = wmask & out; // @[AMOALU.scala 104:19]
  assign _T_93 = ~wmask & io_lhs; // @[AMOALU.scala 104:34]
  assign io_out = _T_91 | _T_93; // @[AMOALU.scala 104:10]
  assign AMOALU_covSum = 30'h0;
  assign io_covSum = AMOALU_covSum;
  assign metaAssert = 1'h0;
endmodule
module ICache(
  input         clock,
  input         reset,
  input         auto_master_out_a_ready,
  output        auto_master_out_a_valid,
  output [31:0] auto_master_out_a_bits_address,
  input         auto_master_out_d_valid,
  input  [2:0]  auto_master_out_d_bits_opcode,
  input  [3:0]  auto_master_out_d_bits_size,
  input  [63:0] auto_master_out_d_bits_data,
  input         auto_master_out_d_bits_corrupt,
  output        io_req_ready,
  input         io_req_valid,
  input  [38:0] io_req_bits_addr,
  input  [31:0] io_s1_paddr,
  input         io_s1_kill,
  input         io_s2_kill,
  output        io_resp_valid,
  output [31:0] io_resp_bits_data,
  output        io_resp_bits_replay,
  output        io_resp_bits_ae,
  input         io_invalidate,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         MaxPeriodFibonacciLFSR_halt
);
  wire  MaxPeriodFibonacciLFSR_clock; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_reset; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_increment; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_0; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_1; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_2; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_3; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_4; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_5; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_6; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_7; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_8; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_9; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_10; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_11; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_12; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_13; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_14; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_15; // @[PRNG.scala 82:22]
  wire [29:0] MaxPeriodFibonacciLFSR_io_covSum; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_metaAssert; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_metaReset; // @[PRNG.scala 82:22]
  reg [20:0] tag_array_0 [0:63]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_0;
  wire [20:0] tag_array_0_tag_rdata_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_0_tag_rdata_addr; // @[DescribedSRAM.scala 23:26]
  wire [20:0] tag_array_0__T_80_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_0__T_80_addr; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_0__T_80_mask; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_0__T_80_en; // @[DescribedSRAM.scala 23:26]
  reg  tag_array_0_tag_rdata_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] tag_array_0_tag_rdata_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg [20:0] tag_array_1 [0:63]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_3;
  wire [20:0] tag_array_1_tag_rdata_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_1_tag_rdata_addr; // @[DescribedSRAM.scala 23:26]
  wire [20:0] tag_array_1__T_80_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_1__T_80_addr; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_1__T_80_mask; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_1__T_80_en; // @[DescribedSRAM.scala 23:26]
  reg  tag_array_1_tag_rdata_en_pipe_0;
  reg [31:0] _RAND_4;
  reg [5:0] tag_array_1_tag_rdata_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [20:0] tag_array_2 [0:63]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_6;
  wire [20:0] tag_array_2_tag_rdata_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_2_tag_rdata_addr; // @[DescribedSRAM.scala 23:26]
  wire [20:0] tag_array_2__T_80_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_2__T_80_addr; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_2__T_80_mask; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_2__T_80_en; // @[DescribedSRAM.scala 23:26]
  reg  tag_array_2_tag_rdata_en_pipe_0;
  reg [31:0] _RAND_7;
  reg [5:0] tag_array_2_tag_rdata_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [20:0] tag_array_3 [0:63]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_9;
  wire [20:0] tag_array_3_tag_rdata_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_3_tag_rdata_addr; // @[DescribedSRAM.scala 23:26]
  wire [20:0] tag_array_3__T_80_data; // @[DescribedSRAM.scala 23:26]
  wire [5:0] tag_array_3__T_80_addr; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_3__T_80_mask; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_3__T_80_en; // @[DescribedSRAM.scala 23:26]
  reg  tag_array_3_tag_rdata_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [5:0] tag_array_3_tag_rdata_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [31:0] data_arrays_0_0 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_12;
  wire [31:0] data_arrays_0_0__T_262_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_0__T_262_addr; // @[DescribedSRAM.scala 23:26]
  wire [31:0] data_arrays_0_0__T_256_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_0__T_256_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_0__T_256_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_0__T_256_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_0__T_262_en_pipe_0;
  reg [31:0] _RAND_13;
  reg [8:0] data_arrays_0_0__T_262_addr_pipe_0;
  reg [31:0] _RAND_14;
  reg [31:0] data_arrays_0_1 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_15;
  wire [31:0] data_arrays_0_1__T_262_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_1__T_262_addr; // @[DescribedSRAM.scala 23:26]
  wire [31:0] data_arrays_0_1__T_256_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_1__T_256_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_1__T_256_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_1__T_256_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_1__T_262_en_pipe_0;
  reg [31:0] _RAND_16;
  reg [8:0] data_arrays_0_1__T_262_addr_pipe_0;
  reg [31:0] _RAND_17;
  reg [31:0] data_arrays_0_2 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_18;
  wire [31:0] data_arrays_0_2__T_262_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_2__T_262_addr; // @[DescribedSRAM.scala 23:26]
  wire [31:0] data_arrays_0_2__T_256_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_2__T_256_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_2__T_256_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_2__T_256_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_2__T_262_en_pipe_0;
  reg [31:0] _RAND_19;
  reg [8:0] data_arrays_0_2__T_262_addr_pipe_0;
  reg [31:0] _RAND_20;
  reg [31:0] data_arrays_0_3 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_21;
  wire [31:0] data_arrays_0_3__T_262_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_3__T_262_addr; // @[DescribedSRAM.scala 23:26]
  wire [31:0] data_arrays_0_3__T_256_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_0_3__T_256_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_3__T_256_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_0_3__T_256_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_0_3__T_262_en_pipe_0;
  reg [31:0] _RAND_22;
  reg [8:0] data_arrays_0_3__T_262_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [31:0] data_arrays_1_0 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_24;
  wire [31:0] data_arrays_1_0__T_300_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_1_0__T_300_addr; // @[DescribedSRAM.scala 23:26]
  wire [31:0] data_arrays_1_0__T_294_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_1_0__T_294_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_1_0__T_294_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_1_0__T_294_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_1_0__T_300_en_pipe_0;
  reg [31:0] _RAND_25;
  reg [8:0] data_arrays_1_0__T_300_addr_pipe_0;
  reg [31:0] _RAND_26;
  reg [31:0] data_arrays_1_1 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_27;
  wire [31:0] data_arrays_1_1__T_300_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_1_1__T_300_addr; // @[DescribedSRAM.scala 23:26]
  wire [31:0] data_arrays_1_1__T_294_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_1_1__T_294_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_1_1__T_294_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_1_1__T_294_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_1_1__T_300_en_pipe_0;
  reg [31:0] _RAND_28;
  reg [8:0] data_arrays_1_1__T_300_addr_pipe_0;
  reg [31:0] _RAND_29;
  reg [31:0] data_arrays_1_2 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_30;
  wire [31:0] data_arrays_1_2__T_300_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_1_2__T_300_addr; // @[DescribedSRAM.scala 23:26]
  wire [31:0] data_arrays_1_2__T_294_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_1_2__T_294_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_1_2__T_294_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_1_2__T_294_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_1_2__T_300_en_pipe_0;
  reg [31:0] _RAND_31;
  reg [8:0] data_arrays_1_2__T_300_addr_pipe_0;
  reg [31:0] _RAND_32;
  reg [31:0] data_arrays_1_3 [0:511]; // @[DescribedSRAM.scala 23:26]
  reg [31:0] _RAND_33;
  wire [31:0] data_arrays_1_3__T_300_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_1_3__T_300_addr; // @[DescribedSRAM.scala 23:26]
  wire [31:0] data_arrays_1_3__T_294_data; // @[DescribedSRAM.scala 23:26]
  wire [8:0] data_arrays_1_3__T_294_addr; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_1_3__T_294_mask; // @[DescribedSRAM.scala 23:26]
  wire  data_arrays_1_3__T_294_en; // @[DescribedSRAM.scala 23:26]
  reg  data_arrays_1_3__T_300_en_pipe_0;
  reg [31:0] _RAND_34;
  reg [8:0] data_arrays_1_3__T_300_addr_pipe_0;
  reg [31:0] _RAND_35;
  wire  s0_valid; // @[Decoupled.scala 40:37]
  reg  s1_valid; // @[ICache.scala 166:21]
  reg [31:0] _RAND_36;
  reg [255:0] vb_array; // @[ICache.scala 228:21]
  reg [255:0] _RAND_37;
  wire [6:0] _T_109; // @[Cat.scala 29:58]
  wire [255:0] _T_110; // @[ICache.scala 256:25]
  wire  _T_116; // @[ICache.scala 259:33]
  wire  s1_tag_hit_0; // @[ICache.scala 259:26]
  wire [6:0] _T_137; // @[Cat.scala 29:58]
  wire [255:0] _T_138; // @[ICache.scala 256:25]
  wire  _T_144; // @[ICache.scala 259:33]
  wire  s1_tag_hit_1; // @[ICache.scala 259:26]
  wire  _T; // @[ICache.scala 169:35]
  wire [7:0] _T_165; // @[Cat.scala 29:58]
  wire [255:0] _T_166; // @[ICache.scala 256:25]
  wire  _T_172; // @[ICache.scala 259:33]
  wire  s1_tag_hit_2; // @[ICache.scala 259:26]
  wire  _T_1; // @[ICache.scala 169:35]
  wire [7:0] _T_193; // @[Cat.scala 29:58]
  wire [255:0] _T_194; // @[ICache.scala 256:25]
  wire  _T_200; // @[ICache.scala 259:33]
  wire  s1_tag_hit_3; // @[ICache.scala 259:26]
  wire  _T_5; // @[ICache.scala 171:35]
  reg  s2_valid; // @[ICache.scala 171:25]
  reg [31:0] _RAND_38;
  reg  s2_hit; // @[ICache.scala 172:23]
  reg [31:0] _RAND_39;
  reg  invalidated; // @[ICache.scala 174:24]
  reg [31:0] _RAND_40;
  reg  refill_valid; // @[ICache.scala 175:29]
  reg [31:0] _RAND_41;
  wire  _T_9; // @[ICache.scala 179:26]
  wire  s2_miss; // @[ICache.scala 179:37]
  reg  _T_12; // @[ICache.scala 181:45]
  reg [31:0] _RAND_42;
  wire  s2_request_refill; // @[ICache.scala 181:35]
  wire  refill_fire; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ICache.scala 180:41]
  wire  s1_can_request_refill; // @[ICache.scala 180:31]
  wire  _T_13; // @[ICache.scala 182:54]
  reg [31:0] refill_paddr; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  wire [19:0] refill_tag; // @[ICache.scala 184:33]
  wire [5:0] refill_idx; // @[ICache.scala 480:21]
  wire  refill_one_beat; // @[ICache.scala 186:41]
  wire [26:0] _T_22; // @[package.scala 212:77]
  wire [8:0] _T_25; // @[Edges.scala 221:59]
  wire [8:0] _T_27; // @[Edges.scala 222:14]
  reg [8:0] _T_28; // @[Edges.scala 230:27]
  reg [31:0] _RAND_44;
  wire [8:0] _T_30; // @[Edges.scala 231:28]
  wire  _T_31; // @[Edges.scala 232:25]
  wire  _T_32; // @[Edges.scala 233:25]
  wire  _T_33; // @[Edges.scala 233:47]
  wire  _T_34; // @[Edges.scala 233:37]
  wire  d_done; // @[Edges.scala 234:22]
  wire [8:0] refill_cnt; // @[Edges.scala 235:25]
  wire  refill_done; // @[ICache.scala 192:37]
  wire [7:0] _T_44; // @[PRNG.scala 86:17]
  wire [15:0] _T_52; // @[PRNG.scala 86:17]
  wire [1:0] repl_way; // @[ICache.scala 198:35]
  wire [7:0] _T_55; // @[Cat.scala 29:58]
  reg  accruedRefillError; // @[ICache.scala 216:31]
  reg [31:0] _RAND_45;
  wire  _T_72; // @[ICache.scala 217:58]
  wire  _T_73; // @[ICache.scala 217:62]
  wire  refillError; // @[ICache.scala 217:43]
  wire  _T_88; // @[ICache.scala 232:72]
  wire [255:0] _T_89; // @[ICache.scala 232:32]
  wire [255:0] _T_90; // @[ICache.scala 232:32]
  wire [255:0] _T_92; // @[ICache.scala 232:32]
  wire  s2_tag_disparity; // @[ICache.scala 305:72]
  wire  _T_338; // @[ICache.scala 328:22]
  wire  invalidate; // @[ICache.scala 328:39]
  wire  _GEN_30; // @[ICache.scala 235:21]
  wire  s1_tl_error_0; // @[ICache.scala 261:32]
  wire  s1_tl_error_1; // @[ICache.scala 261:32]
  wire  s1_tl_error_2; // @[ICache.scala 261:32]
  wire  s1_tl_error_3; // @[ICache.scala 261:32]
  wire [1:0] _T_217; // @[Bitwise.scala 47:55]
  wire [1:0] _T_219; // @[Bitwise.scala 47:55]
  wire [2:0] _T_221; // @[Bitwise.scala 47:55]
  wire  _T_223; // @[ICache.scala 264:115]
  wire  _T_224; // @[ICache.scala 264:39]
  wire  _T_226; // @[ICache.scala 264:9]
  wire  _T_230; // @[ICache.scala 281:28]
  wire  _T_235; // @[ICache.scala 282:32]
  wire [8:0] _T_240; // @[ICache.scala 283:52]
  wire [8:0] _T_241; // @[ICache.scala 283:79]
  wire [31:0] _GEN_54; // @[ICache.scala 293:71]
  wire [31:0] _GEN_55; // @[ICache.scala 293:71]
  wire [31:0] _GEN_56; // @[ICache.scala 293:71]
  wire [31:0] _GEN_57; // @[ICache.scala 293:71]
  wire  _T_268; // @[ICache.scala 281:28]
  reg  s2_tag_hit_0; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg  s2_tag_hit_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg  s2_tag_hit_2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg  s2_tag_hit_3; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [31:0] s2_dout_0; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [31:0] s2_dout_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [31:0] s2_dout_2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [31:0] s2_dout_3; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  wire [31:0] _T_315; // @[Mux.scala 27:72]
  wire [31:0] _T_316; // @[Mux.scala 27:72]
  wire [31:0] _T_317; // @[Mux.scala 27:72]
  wire [31:0] _T_318; // @[Mux.scala 27:72]
  wire [31:0] _T_319; // @[Mux.scala 27:72]
  wire [31:0] _T_320; // @[Mux.scala 27:72]
  wire [3:0] _T_328; // @[ICache.scala 306:43]
  wire  _T_329; // @[ICache.scala 306:50]
  reg  s2_tl_error; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  wire  _GEN_101; // @[ICache.scala 471:22]
  reg [5:0] ICache_state; // @[Register tracking ICache state]
  reg [31:0] _RAND_55;
  reg  ICache_cov [0:63]; // @[Coverage map for ICache]
  reg [31:0] _RAND_56;
  wire  ICache_cov_read_data; // @[Coverage map for ICache]
  wire [5:0] ICache_cov_read_addr; // @[Coverage map for ICache]
  wire  ICache_cov_write_data; // @[Coverage map for ICache]
  wire [5:0] ICache_cov_write_addr; // @[Coverage map for ICache]
  wire  ICache_cov_write_mask; // @[Coverage map for ICache]
  wire  ICache_cov_write_en; // @[Coverage map for ICache]
  reg [29:0] ICache_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_57;
  wire  s2_hit_shl;
  wire [5:0] s2_hit_pad;
  wire [1:0] s2_valid_shl;
  wire [5:0] s2_valid_pad;
  wire [2:0] refill_valid_shl;
  wire [5:0] refill_valid_pad;
  wire [3:0] s1_valid_shl;
  wire [5:0] s1_valid_pad;
  wire [4:0] invalidated_shl;
  wire [5:0] invalidated_pad;
  wire [5:0] s2_tag_hit_0_shl;
  wire [5:0] s2_tag_hit_0_pad;
  wire [5:0] s2_tag_hit_1_shl;
  wire [5:0] s2_tag_hit_1_pad;
  wire [5:0] s2_tag_hit_2_shl;
  wire [5:0] s2_tag_hit_2_pad;
  wire [5:0] s2_tag_hit_3_shl;
  wire [5:0] s2_tag_hit_3_pad;
  wire [5:0] ICache_xor3;
  wire [5:0] ICache_xor4;
  wire [5:0] ICache_xor1;
  wire [5:0] ICache_xor5;
  wire [5:0] ICache_xor14;
  wire [5:0] ICache_xor6;
  wire [5:0] ICache_xor2;
  wire [5:0] ICache_xor0;
  wire [29:0] MaxPeriodFibonacciLFSR_sum;
  wire  stopEn0;
  wire  MaxPeriodFibonacciLFSR_metaAssert_wire;
  wire  ICache_or0;
  reg  ICache_metaAssert;
  reg [31:0] _RAND_58;
  MaxPeriodFibonacciLFSR MaxPeriodFibonacciLFSR ( // @[PRNG.scala 82:22]
    .clock(MaxPeriodFibonacciLFSR_clock),
    .reset(MaxPeriodFibonacciLFSR_reset),
    .io_increment(MaxPeriodFibonacciLFSR_io_increment),
    .io_out_0(MaxPeriodFibonacciLFSR_io_out_0),
    .io_out_1(MaxPeriodFibonacciLFSR_io_out_1),
    .io_out_2(MaxPeriodFibonacciLFSR_io_out_2),
    .io_out_3(MaxPeriodFibonacciLFSR_io_out_3),
    .io_out_4(MaxPeriodFibonacciLFSR_io_out_4),
    .io_out_5(MaxPeriodFibonacciLFSR_io_out_5),
    .io_out_6(MaxPeriodFibonacciLFSR_io_out_6),
    .io_out_7(MaxPeriodFibonacciLFSR_io_out_7),
    .io_out_8(MaxPeriodFibonacciLFSR_io_out_8),
    .io_out_9(MaxPeriodFibonacciLFSR_io_out_9),
    .io_out_10(MaxPeriodFibonacciLFSR_io_out_10),
    .io_out_11(MaxPeriodFibonacciLFSR_io_out_11),
    .io_out_12(MaxPeriodFibonacciLFSR_io_out_12),
    .io_out_13(MaxPeriodFibonacciLFSR_io_out_13),
    .io_out_14(MaxPeriodFibonacciLFSR_io_out_14),
    .io_out_15(MaxPeriodFibonacciLFSR_io_out_15),
    .io_covSum(MaxPeriodFibonacciLFSR_io_covSum),
    .metaAssert(MaxPeriodFibonacciLFSR_metaAssert),
    .metaReset(MaxPeriodFibonacciLFSR_metaReset)
  );
  assign tag_array_0_tag_rdata_addr = tag_array_0_tag_rdata_addr_pipe_0;
  assign tag_array_0_tag_rdata_data = tag_array_0[tag_array_0_tag_rdata_addr]; // @[DescribedSRAM.scala 23:26]
  assign tag_array_0__T_80_data = {refillError,refill_tag};
  assign tag_array_0__T_80_addr = refill_paddr[11:6];
  assign tag_array_0__T_80_mask = repl_way == 2'h0;
  assign tag_array_0__T_80_en = refill_one_beat & d_done;
  assign tag_array_1_tag_rdata_addr = tag_array_1_tag_rdata_addr_pipe_0;
  assign tag_array_1_tag_rdata_data = tag_array_1[tag_array_1_tag_rdata_addr]; // @[DescribedSRAM.scala 23:26]
  assign tag_array_1__T_80_data = {refillError,refill_tag};
  assign tag_array_1__T_80_addr = refill_paddr[11:6];
  assign tag_array_1__T_80_mask = repl_way == 2'h1;
  assign tag_array_1__T_80_en = refill_one_beat & d_done;
  assign tag_array_2_tag_rdata_addr = tag_array_2_tag_rdata_addr_pipe_0;
  assign tag_array_2_tag_rdata_data = tag_array_2[tag_array_2_tag_rdata_addr]; // @[DescribedSRAM.scala 23:26]
  assign tag_array_2__T_80_data = {refillError,refill_tag};
  assign tag_array_2__T_80_addr = refill_paddr[11:6];
  assign tag_array_2__T_80_mask = repl_way == 2'h2;
  assign tag_array_2__T_80_en = refill_one_beat & d_done;
  assign tag_array_3_tag_rdata_addr = tag_array_3_tag_rdata_addr_pipe_0;
  assign tag_array_3_tag_rdata_data = tag_array_3[tag_array_3_tag_rdata_addr]; // @[DescribedSRAM.scala 23:26]
  assign tag_array_3__T_80_data = {refillError,refill_tag};
  assign tag_array_3__T_80_addr = refill_paddr[11:6];
  assign tag_array_3__T_80_mask = repl_way == 2'h3;
  assign tag_array_3__T_80_en = refill_one_beat & d_done;
  assign data_arrays_0_0__T_262_addr = data_arrays_0_0__T_262_addr_pipe_0;
  assign data_arrays_0_0__T_262_data = data_arrays_0_0[data_arrays_0_0__T_262_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_0__T_256_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_0__T_256_addr = refill_one_beat ? _T_241 : io_req_bits_addr[11:3];
  assign data_arrays_0_0__T_256_mask = repl_way == 2'h0;
  assign data_arrays_0_0__T_256_en = refill_one_beat & ~invalidated;
  assign data_arrays_0_1__T_262_addr = data_arrays_0_1__T_262_addr_pipe_0;
  assign data_arrays_0_1__T_262_data = data_arrays_0_1[data_arrays_0_1__T_262_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_1__T_256_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_1__T_256_addr = refill_one_beat ? _T_241 : io_req_bits_addr[11:3];
  assign data_arrays_0_1__T_256_mask = repl_way == 2'h1;
  assign data_arrays_0_1__T_256_en = refill_one_beat & ~invalidated;
  assign data_arrays_0_2__T_262_addr = data_arrays_0_2__T_262_addr_pipe_0;
  assign data_arrays_0_2__T_262_data = data_arrays_0_2[data_arrays_0_2__T_262_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_2__T_256_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_2__T_256_addr = refill_one_beat ? _T_241 : io_req_bits_addr[11:3];
  assign data_arrays_0_2__T_256_mask = repl_way == 2'h2;
  assign data_arrays_0_2__T_256_en = refill_one_beat & ~invalidated;
  assign data_arrays_0_3__T_262_addr = data_arrays_0_3__T_262_addr_pipe_0;
  assign data_arrays_0_3__T_262_data = data_arrays_0_3[data_arrays_0_3__T_262_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_0_3__T_256_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_3__T_256_addr = refill_one_beat ? _T_241 : io_req_bits_addr[11:3];
  assign data_arrays_0_3__T_256_mask = repl_way == 2'h3;
  assign data_arrays_0_3__T_256_en = refill_one_beat & ~invalidated;
  assign data_arrays_1_0__T_300_addr = data_arrays_1_0__T_300_addr_pipe_0;
  assign data_arrays_1_0__T_300_data = data_arrays_1_0[data_arrays_1_0__T_300_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_1_0__T_294_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_0__T_294_addr = refill_one_beat ? _T_241 : io_req_bits_addr[11:3];
  assign data_arrays_1_0__T_294_mask = repl_way == 2'h0;
  assign data_arrays_1_0__T_294_en = refill_one_beat & ~invalidated;
  assign data_arrays_1_1__T_300_addr = data_arrays_1_1__T_300_addr_pipe_0;
  assign data_arrays_1_1__T_300_data = data_arrays_1_1[data_arrays_1_1__T_300_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_1_1__T_294_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_1__T_294_addr = refill_one_beat ? _T_241 : io_req_bits_addr[11:3];
  assign data_arrays_1_1__T_294_mask = repl_way == 2'h1;
  assign data_arrays_1_1__T_294_en = refill_one_beat & ~invalidated;
  assign data_arrays_1_2__T_300_addr = data_arrays_1_2__T_300_addr_pipe_0;
  assign data_arrays_1_2__T_300_data = data_arrays_1_2[data_arrays_1_2__T_300_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_1_2__T_294_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_2__T_294_addr = refill_one_beat ? _T_241 : io_req_bits_addr[11:3];
  assign data_arrays_1_2__T_294_mask = repl_way == 2'h2;
  assign data_arrays_1_2__T_294_en = refill_one_beat & ~invalidated;
  assign data_arrays_1_3__T_300_addr = data_arrays_1_3__T_300_addr_pipe_0;
  assign data_arrays_1_3__T_300_data = data_arrays_1_3[data_arrays_1_3__T_300_addr]; // @[DescribedSRAM.scala 23:26]
  assign data_arrays_1_3__T_294_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_3__T_294_addr = refill_one_beat ? _T_241 : io_req_bits_addr[11:3];
  assign data_arrays_1_3__T_294_mask = repl_way == 2'h3;
  assign data_arrays_1_3__T_294_en = refill_one_beat & ~invalidated;
  assign s0_valid = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37]
  assign _T_109 = {1'h0,io_s1_paddr[11:6]}; // @[Cat.scala 29:58]
  assign _T_110 = vb_array >> _T_109; // @[ICache.scala 256:25]
  assign _T_116 = tag_array_0_tag_rdata_data[19:0] == io_s1_paddr[31:12]; // @[ICache.scala 259:33]
  assign s1_tag_hit_0 = _T_110[0] & _T_116; // @[ICache.scala 259:26]
  assign _T_137 = {1'h1,io_s1_paddr[11:6]}; // @[Cat.scala 29:58]
  assign _T_138 = vb_array >> _T_137; // @[ICache.scala 256:25]
  assign _T_144 = tag_array_1_tag_rdata_data[19:0] == io_s1_paddr[31:12]; // @[ICache.scala 259:33]
  assign s1_tag_hit_1 = _T_138[0] & _T_144; // @[ICache.scala 259:26]
  assign _T = s1_tag_hit_0 | s1_tag_hit_1; // @[ICache.scala 169:35]
  assign _T_165 = {2'h2,io_s1_paddr[11:6]}; // @[Cat.scala 29:58]
  assign _T_166 = vb_array >> _T_165; // @[ICache.scala 256:25]
  assign _T_172 = tag_array_2_tag_rdata_data[19:0] == io_s1_paddr[31:12]; // @[ICache.scala 259:33]
  assign s1_tag_hit_2 = _T_166[0] & _T_172; // @[ICache.scala 259:26]
  assign _T_1 = _T | s1_tag_hit_2; // @[ICache.scala 169:35]
  assign _T_193 = {2'h3,io_s1_paddr[11:6]}; // @[Cat.scala 29:58]
  assign _T_194 = vb_array >> _T_193; // @[ICache.scala 256:25]
  assign _T_200 = tag_array_3_tag_rdata_data[19:0] == io_s1_paddr[31:12]; // @[ICache.scala 259:33]
  assign s1_tag_hit_3 = _T_194[0] & _T_200; // @[ICache.scala 259:26]
  assign _T_5 = s1_valid & ~io_s1_kill; // @[ICache.scala 171:35]
  assign _T_9 = s2_valid & ~s2_hit; // @[ICache.scala 179:26]
  assign s2_miss = _T_9 & ~io_s2_kill; // @[ICache.scala 179:37]
  assign s2_request_refill = s2_miss & _T_12; // @[ICache.scala 181:35]
  assign refill_fire = auto_master_out_a_ready & s2_request_refill; // @[Decoupled.scala 40:37]
  assign _T_11 = s2_miss | refill_valid; // @[ICache.scala 180:41]
  assign s1_can_request_refill = ~_T_11; // @[ICache.scala 180:31]
  assign _T_13 = s1_valid & s1_can_request_refill; // @[ICache.scala 182:54]
  assign refill_tag = refill_paddr[31:12]; // @[ICache.scala 184:33]
  assign refill_idx = refill_paddr[11:6]; // @[ICache.scala 480:21]
  assign refill_one_beat = auto_master_out_d_valid & auto_master_out_d_bits_opcode[0]; // @[ICache.scala 186:41]
  assign _T_22 = 27'hfff << auto_master_out_d_bits_size; // @[package.scala 212:77]
  assign _T_25 = ~_T_22[11:3]; // @[Edges.scala 221:59]
  assign _T_27 = auto_master_out_d_bits_opcode[0] ? _T_25 : 9'h0; // @[Edges.scala 222:14]
  assign _T_30 = _T_28 - 9'h1; // @[Edges.scala 231:28]
  assign _T_31 = _T_28 == 9'h0; // @[Edges.scala 232:25]
  assign _T_32 = _T_28 == 9'h1; // @[Edges.scala 233:25]
  assign _T_33 = _T_27 == 9'h0; // @[Edges.scala 233:47]
  assign _T_34 = _T_32 | _T_33; // @[Edges.scala 233:37]
  assign d_done = _T_34 & auto_master_out_d_valid; // @[Edges.scala 234:22]
  assign refill_cnt = _T_27 & ~_T_30; // @[Edges.scala 235:25]
  assign refill_done = refill_one_beat & d_done; // @[ICache.scala 192:37]
  assign _T_44 = {MaxPeriodFibonacciLFSR_io_out_7,MaxPeriodFibonacciLFSR_io_out_6,MaxPeriodFibonacciLFSR_io_out_5,MaxPeriodFibonacciLFSR_io_out_4,MaxPeriodFibonacciLFSR_io_out_3,MaxPeriodFibonacciLFSR_io_out_2,MaxPeriodFibonacciLFSR_io_out_1,MaxPeriodFibonacciLFSR_io_out_0}; // @[PRNG.scala 86:17]
  assign _T_52 = {MaxPeriodFibonacciLFSR_io_out_15,MaxPeriodFibonacciLFSR_io_out_14,MaxPeriodFibonacciLFSR_io_out_13,MaxPeriodFibonacciLFSR_io_out_12,MaxPeriodFibonacciLFSR_io_out_11,MaxPeriodFibonacciLFSR_io_out_10,MaxPeriodFibonacciLFSR_io_out_9,MaxPeriodFibonacciLFSR_io_out_8,_T_44}; // @[PRNG.scala 86:17]
  assign repl_way = _T_52[1:0]; // @[ICache.scala 198:35]
  assign _T_55 = {repl_way,refill_idx}; // @[Cat.scala 29:58]
  assign _T_72 = refill_cnt > 9'h0; // @[ICache.scala 217:58]
  assign _T_73 = _T_72 & accruedRefillError; // @[ICache.scala 217:62]
  assign refillError = auto_master_out_d_bits_corrupt | _T_73; // @[ICache.scala 217:43]
  assign _T_88 = refill_done & ~invalidated; // @[ICache.scala 232:72]
  assign _T_89 = 256'h1 << _T_55; // @[ICache.scala 232:32]
  assign _T_90 = vb_array | _T_89; // @[ICache.scala 232:32]
  assign _T_92 = ~vb_array | _T_89; // @[ICache.scala 232:32]
  assign s2_tag_disparity = |4'h0; // @[ICache.scala 305:72]
  assign _T_338 = s2_valid & s2_tag_disparity; // @[ICache.scala 328:22]
  assign invalidate = _T_338 | io_invalidate; // @[ICache.scala 328:39]
  assign _GEN_30 = invalidate | invalidated; // @[ICache.scala 235:21]
  assign s1_tl_error_0 = s1_tag_hit_0 & tag_array_0_tag_rdata_data[20]; // @[ICache.scala 261:32]
  assign s1_tl_error_1 = s1_tag_hit_1 & tag_array_1_tag_rdata_data[20]; // @[ICache.scala 261:32]
  assign s1_tl_error_2 = s1_tag_hit_2 & tag_array_2_tag_rdata_data[20]; // @[ICache.scala 261:32]
  assign s1_tl_error_3 = s1_tag_hit_3 & tag_array_3_tag_rdata_data[20]; // @[ICache.scala 261:32]
  assign _T_217 = s1_tag_hit_0 + s1_tag_hit_1; // @[Bitwise.scala 47:55]
  assign _T_219 = s1_tag_hit_2 + s1_tag_hit_3; // @[Bitwise.scala 47:55]
  assign _T_221 = _T_217 + _T_219; // @[Bitwise.scala 47:55]
  assign _T_223 = _T_221 <= 3'h1; // @[ICache.scala 264:115]
  assign _T_224 = ~s1_valid | _T_223; // @[ICache.scala 264:39]
  assign _T_226 = _T_224 | reset; // @[ICache.scala 264:9]
  assign _T_230 = s0_valid & ~io_req_bits_addr[2]; // @[ICache.scala 281:28]
  assign _T_235 = refill_one_beat & ~invalidated; // @[ICache.scala 282:32]
  assign _T_240 = {refill_idx, 3'h0}; // @[ICache.scala 283:52]
  assign _T_241 = _T_240 | refill_cnt; // @[ICache.scala 283:79]
  assign _GEN_54 = data_arrays_0_0__T_262_data; // @[ICache.scala 293:71]
  assign _GEN_55 = data_arrays_0_1__T_262_data; // @[ICache.scala 293:71]
  assign _GEN_56 = data_arrays_0_2__T_262_data; // @[ICache.scala 293:71]
  assign _GEN_57 = data_arrays_0_3__T_262_data; // @[ICache.scala 293:71]
  assign _T_268 = s0_valid & io_req_bits_addr[2]; // @[ICache.scala 281:28]
  assign _T_315 = s2_tag_hit_0 ? s2_dout_0 : 32'h0; // @[Mux.scala 27:72]
  assign _T_316 = s2_tag_hit_1 ? s2_dout_1 : 32'h0; // @[Mux.scala 27:72]
  assign _T_317 = s2_tag_hit_2 ? s2_dout_2 : 32'h0; // @[Mux.scala 27:72]
  assign _T_318 = s2_tag_hit_3 ? s2_dout_3 : 32'h0; // @[Mux.scala 27:72]
  assign _T_319 = _T_315 | _T_316; // @[Mux.scala 27:72]
  assign _T_320 = _T_319 | _T_317; // @[Mux.scala 27:72]
  assign _T_328 = {s1_tl_error_3,s1_tl_error_2,s1_tl_error_1,s1_tl_error_0}; // @[ICache.scala 306:43]
  assign _T_329 = |_T_328; // @[ICache.scala 306:50]
  assign _GEN_101 = refill_fire | refill_valid; // @[ICache.scala 471:22]
  assign auto_master_out_a_valid = s2_miss & _T_12; // @[LazyModule.scala 305:12]
  assign auto_master_out_a_bits_address = {refill_paddr[31:6], 6'h0}; // @[LazyModule.scala 305:12]
  assign io_req_ready = ~refill_one_beat; // @[ICache.scala 188:16]
  assign io_resp_valid = s2_valid & s2_hit; // @[ICache.scala 333:21]
  assign io_resp_bits_data = _T_320 | _T_318; // @[ICache.scala 330:25]
  assign io_resp_bits_replay = |4'h0; // @[ICache.scala 332:27]
  assign io_resp_bits_ae = s2_tl_error; // @[ICache.scala 331:23]
  assign MaxPeriodFibonacciLFSR_clock = clock;
  assign MaxPeriodFibonacciLFSR_reset = reset;
  assign MaxPeriodFibonacciLFSR_io_increment = auto_master_out_a_ready & s2_request_refill; // @[PRNG.scala 85:23]
  assign ICache_cov_read_addr = ICache_state;
  assign ICache_cov_read_data = ICache_cov[ICache_cov_read_addr]; // @[Coverage map for ICache]
  assign ICache_cov_write_data = 1'h1;
  assign ICache_cov_write_addr = ICache_state;
  assign ICache_cov_write_mask = 1'h1;
  assign ICache_cov_write_en = 1'h1;
  assign s2_hit_shl = s2_hit;
  assign s2_hit_pad = {5'h0,s2_hit_shl};
  assign s2_valid_shl = {s2_valid, 1'h0};
  assign s2_valid_pad = {4'h0,s2_valid_shl};
  assign refill_valid_shl = {refill_valid, 2'h0};
  assign refill_valid_pad = {3'h0,refill_valid_shl};
  assign s1_valid_shl = {s1_valid, 3'h0};
  assign s1_valid_pad = {2'h0,s1_valid_shl};
  assign invalidated_shl = {invalidated, 4'h0};
  assign invalidated_pad = {1'h0,invalidated_shl};
  assign s2_tag_hit_0_shl = {s2_tag_hit_0, 5'h0};
  assign s2_tag_hit_0_pad = s2_tag_hit_0_shl;
  assign s2_tag_hit_1_shl = {s2_tag_hit_1, 5'h0};
  assign s2_tag_hit_1_pad = s2_tag_hit_1_shl;
  assign s2_tag_hit_2_shl = {s2_tag_hit_2, 5'h0};
  assign s2_tag_hit_2_pad = s2_tag_hit_2_shl;
  assign s2_tag_hit_3_shl = {s2_tag_hit_3, 5'h0};
  assign s2_tag_hit_3_pad = s2_tag_hit_3_shl;
  assign ICache_xor3 = s2_hit_pad ^ s2_valid_pad;
  assign ICache_xor4 = refill_valid_pad ^ s1_valid_pad;
  assign ICache_xor1 = ICache_xor3 ^ ICache_xor4;
  assign ICache_xor5 = invalidated_pad ^ s2_tag_hit_0_pad;
  assign ICache_xor14 = s2_tag_hit_2_pad ^ s2_tag_hit_3_pad;
  assign ICache_xor6 = s2_tag_hit_1_pad ^ ICache_xor14;
  assign ICache_xor2 = ICache_xor5 ^ ICache_xor6;
  assign ICache_xor0 = ICache_xor1 ^ ICache_xor2;
  assign MaxPeriodFibonacciLFSR_sum = ICache_covSum + MaxPeriodFibonacciLFSR_io_covSum;
  assign io_covSum = MaxPeriodFibonacciLFSR_sum;
  assign stopEn0 = ~_T_226;
  assign MaxPeriodFibonacciLFSR_metaAssert_wire = MaxPeriodFibonacciLFSR_metaAssert;
  assign ICache_or0 = stopEn0 | MaxPeriodFibonacciLFSR_metaAssert_wire;
  assign metaAssert = ICache_metaAssert;
  assign MaxPeriodFibonacciLFSR_metaReset = metaReset | MaxPeriodFibonacciLFSR_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_0[initvar] = _RAND_0[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tag_array_0_tag_rdata_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tag_array_0_tag_rdata_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_1[initvar] = _RAND_3[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  tag_array_1_tag_rdata_en_pipe_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  tag_array_1_tag_rdata_addr_pipe_0 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_2[initvar] = _RAND_6[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  tag_array_2_tag_rdata_en_pipe_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tag_array_2_tag_rdata_addr_pipe_0 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_3[initvar] = _RAND_9[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  tag_array_3_tag_rdata_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  tag_array_3_tag_rdata_addr_pipe_0 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_0[initvar] = _RAND_12[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  data_arrays_0_0__T_262_en_pipe_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  data_arrays_0_0__T_262_addr_pipe_0 = _RAND_14[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_1[initvar] = _RAND_15[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  data_arrays_0_1__T_262_en_pipe_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  data_arrays_0_1__T_262_addr_pipe_0 = _RAND_17[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_2[initvar] = _RAND_18[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  data_arrays_0_2__T_262_en_pipe_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  data_arrays_0_2__T_262_addr_pipe_0 = _RAND_20[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_3[initvar] = _RAND_21[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  data_arrays_0_3__T_262_en_pipe_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  data_arrays_0_3__T_262_addr_pipe_0 = _RAND_23[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_1_0[initvar] = _RAND_24[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  data_arrays_1_0__T_300_en_pipe_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  data_arrays_1_0__T_300_addr_pipe_0 = _RAND_26[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_1_1[initvar] = _RAND_27[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  data_arrays_1_1__T_300_en_pipe_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  data_arrays_1_1__T_300_addr_pipe_0 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_1_2[initvar] = _RAND_30[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  data_arrays_1_2__T_300_en_pipe_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  data_arrays_1_2__T_300_addr_pipe_0 = _RAND_32[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_1_3[initvar] = _RAND_33[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  data_arrays_1_3__T_300_en_pipe_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  data_arrays_1_3__T_300_addr_pipe_0 = _RAND_35[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  s1_valid = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {8{`RANDOM}};
  vb_array = _RAND_37[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  s2_valid = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  s2_hit = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  invalidated = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  refill_valid = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_12 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  refill_paddr = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_28 = _RAND_44[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  accruedRefillError = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  s2_tag_hit_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  s2_tag_hit_1 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  s2_tag_hit_2 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  s2_tag_hit_3 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  s2_dout_0 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  s2_dout_1 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  s2_dout_2 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  s2_dout_3 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  s2_tl_error = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  ICache_state = _RAND_55[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ICache_cov[initvar] = _RAND_56[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  ICache_covSum = _RAND_57[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  ICache_metaAssert = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(tag_array_0__T_80_en & tag_array_0__T_80_mask) begin
      tag_array_0[tag_array_0__T_80_addr] <= tag_array_0__T_80_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      tag_array_0_tag_rdata_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_0_tag_rdata_en_pipe_0 <= ~refill_done & s0_valid;
    end
    if (metaReset) begin
      tag_array_0_tag_rdata_addr_pipe_0 <= 6'h0;
    end else if (~refill_done & s0_valid) begin
      tag_array_0_tag_rdata_addr_pipe_0 <= io_req_bits_addr[11:6];
    end
    if(tag_array_1__T_80_en & tag_array_1__T_80_mask) begin
      tag_array_1[tag_array_1__T_80_addr] <= tag_array_1__T_80_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      tag_array_1_tag_rdata_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_1_tag_rdata_en_pipe_0 <= ~refill_done & s0_valid;
    end
    if (metaReset) begin
      tag_array_1_tag_rdata_addr_pipe_0 <= 6'h0;
    end else if (~refill_done & s0_valid) begin
      tag_array_1_tag_rdata_addr_pipe_0 <= io_req_bits_addr[11:6];
    end
    if(tag_array_2__T_80_en & tag_array_2__T_80_mask) begin
      tag_array_2[tag_array_2__T_80_addr] <= tag_array_2__T_80_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      tag_array_2_tag_rdata_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_2_tag_rdata_en_pipe_0 <= ~refill_done & s0_valid;
    end
    if (metaReset) begin
      tag_array_2_tag_rdata_addr_pipe_0 <= 6'h0;
    end else if (~refill_done & s0_valid) begin
      tag_array_2_tag_rdata_addr_pipe_0 <= io_req_bits_addr[11:6];
    end
    if(tag_array_3__T_80_en & tag_array_3__T_80_mask) begin
      tag_array_3[tag_array_3__T_80_addr] <= tag_array_3__T_80_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      tag_array_3_tag_rdata_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_3_tag_rdata_en_pipe_0 <= ~refill_done & s0_valid;
    end
    if (metaReset) begin
      tag_array_3_tag_rdata_addr_pipe_0 <= 6'h0;
    end else if (~refill_done & s0_valid) begin
      tag_array_3_tag_rdata_addr_pipe_0 <= io_req_bits_addr[11:6];
    end
    if(data_arrays_0_0__T_256_en & data_arrays_0_0__T_256_mask) begin
      data_arrays_0_0[data_arrays_0_0__T_256_addr] <= data_arrays_0_0__T_256_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_0__T_262_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_0__T_262_en_pipe_0 <= ~_T_235 & _T_230;
    end
    if (metaReset) begin
      data_arrays_0_0__T_262_addr_pipe_0 <= 9'h0;
    end else if (~_T_235 & _T_230) begin
      if (refill_one_beat) begin
        data_arrays_0_0__T_262_addr_pipe_0 <= _T_241;
      end else begin
        data_arrays_0_0__T_262_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_0_1__T_256_en & data_arrays_0_1__T_256_mask) begin
      data_arrays_0_1[data_arrays_0_1__T_256_addr] <= data_arrays_0_1__T_256_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_1__T_262_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_1__T_262_en_pipe_0 <= ~_T_235 & _T_230;
    end
    if (metaReset) begin
      data_arrays_0_1__T_262_addr_pipe_0 <= 9'h0;
    end else if (~_T_235 & _T_230) begin
      if (refill_one_beat) begin
        data_arrays_0_1__T_262_addr_pipe_0 <= _T_241;
      end else begin
        data_arrays_0_1__T_262_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_0_2__T_256_en & data_arrays_0_2__T_256_mask) begin
      data_arrays_0_2[data_arrays_0_2__T_256_addr] <= data_arrays_0_2__T_256_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_2__T_262_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_2__T_262_en_pipe_0 <= ~_T_235 & _T_230;
    end
    if (metaReset) begin
      data_arrays_0_2__T_262_addr_pipe_0 <= 9'h0;
    end else if (~_T_235 & _T_230) begin
      if (refill_one_beat) begin
        data_arrays_0_2__T_262_addr_pipe_0 <= _T_241;
      end else begin
        data_arrays_0_2__T_262_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_0_3__T_256_en & data_arrays_0_3__T_256_mask) begin
      data_arrays_0_3[data_arrays_0_3__T_256_addr] <= data_arrays_0_3__T_256_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_0_3__T_262_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_3__T_262_en_pipe_0 <= ~_T_235 & _T_230;
    end
    if (metaReset) begin
      data_arrays_0_3__T_262_addr_pipe_0 <= 9'h0;
    end else if (~_T_235 & _T_230) begin
      if (refill_one_beat) begin
        data_arrays_0_3__T_262_addr_pipe_0 <= _T_241;
      end else begin
        data_arrays_0_3__T_262_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_1_0__T_294_en & data_arrays_1_0__T_294_mask) begin
      data_arrays_1_0[data_arrays_1_0__T_294_addr] <= data_arrays_1_0__T_294_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_1_0__T_300_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_1_0__T_300_en_pipe_0 <= ~_T_235 & _T_268;
    end
    if (metaReset) begin
      data_arrays_1_0__T_300_addr_pipe_0 <= 9'h0;
    end else if (~_T_235 & _T_268) begin
      if (refill_one_beat) begin
        data_arrays_1_0__T_300_addr_pipe_0 <= _T_241;
      end else begin
        data_arrays_1_0__T_300_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_1_1__T_294_en & data_arrays_1_1__T_294_mask) begin
      data_arrays_1_1[data_arrays_1_1__T_294_addr] <= data_arrays_1_1__T_294_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_1_1__T_300_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_1_1__T_300_en_pipe_0 <= ~_T_235 & _T_268;
    end
    if (metaReset) begin
      data_arrays_1_1__T_300_addr_pipe_0 <= 9'h0;
    end else if (~_T_235 & _T_268) begin
      if (refill_one_beat) begin
        data_arrays_1_1__T_300_addr_pipe_0 <= _T_241;
      end else begin
        data_arrays_1_1__T_300_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_1_2__T_294_en & data_arrays_1_2__T_294_mask) begin
      data_arrays_1_2[data_arrays_1_2__T_294_addr] <= data_arrays_1_2__T_294_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_1_2__T_300_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_1_2__T_300_en_pipe_0 <= ~_T_235 & _T_268;
    end
    if (metaReset) begin
      data_arrays_1_2__T_300_addr_pipe_0 <= 9'h0;
    end else if (~_T_235 & _T_268) begin
      if (refill_one_beat) begin
        data_arrays_1_2__T_300_addr_pipe_0 <= _T_241;
      end else begin
        data_arrays_1_2__T_300_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_1_3__T_294_en & data_arrays_1_3__T_294_mask) begin
      data_arrays_1_3[data_arrays_1_3__T_294_addr] <= data_arrays_1_3__T_294_data; // @[DescribedSRAM.scala 23:26]
    end
    if (metaReset) begin
      data_arrays_1_3__T_300_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_1_3__T_300_en_pipe_0 <= ~_T_235 & _T_268;
    end
    if (metaReset) begin
      data_arrays_1_3__T_300_addr_pipe_0 <= 9'h0;
    end else if (~_T_235 & _T_268) begin
      if (refill_one_beat) begin
        data_arrays_1_3__T_300_addr_pipe_0 <= _T_241;
      end else begin
        data_arrays_1_3__T_300_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if (metaReset) begin
      s1_valid <= 1'h0;
    end else if (reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= s0_valid;
    end
    if (metaReset) begin
      vb_array <= 256'h0;
    end else if (reset) begin
      vb_array <= 256'h0;
    end else if (invalidate) begin
      vb_array <= 256'h0;
    end else if (refill_one_beat) begin
      if (_T_88) begin
        vb_array <= _T_90;
      end else begin
        vb_array <= ~_T_92;
      end
    end
    if (metaReset) begin
      s2_valid <= 1'h0;
    end else if (reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= _T_5;
    end
    if (metaReset) begin
      s2_hit <= 1'h0;
    end else begin
      s2_hit <= _T_1 | s1_tag_hit_3;
    end
    if (metaReset) begin
      invalidated <= 1'h0;
    end else if (~refill_valid) begin
      invalidated <= 1'h0;
    end else begin
      invalidated <= _GEN_30;
    end
    if (metaReset) begin
      refill_valid <= 1'h0;
    end else if (reset) begin
      refill_valid <= 1'h0;
    end else if (refill_done) begin
      refill_valid <= 1'h0;
    end else begin
      refill_valid <= _GEN_101;
    end
    if (metaReset) begin
      _T_12 <= 1'h0;
    end else begin
      _T_12 <= ~_T_11;
    end
    if (metaReset) begin
      refill_paddr <= 32'h0;
    end else if (_T_13) begin
      refill_paddr <= io_s1_paddr;
    end
    if (metaReset) begin
      _T_28 <= 9'h0;
    end else if (reset) begin
      _T_28 <= 9'h0;
    end else if (auto_master_out_d_valid) begin
      if (_T_31) begin
        if (auto_master_out_d_bits_opcode[0]) begin
          _T_28 <= _T_25;
        end else begin
          _T_28 <= 9'h0;
        end
      end else begin
        _T_28 <= _T_30;
      end
    end
    if (metaReset) begin
      accruedRefillError <= 1'h0;
    end else if (refill_one_beat) begin
      accruedRefillError <= refillError;
    end
    if (metaReset) begin
      s2_tag_hit_0 <= 1'h0;
    end else if (s1_valid) begin
      s2_tag_hit_0 <= s1_tag_hit_0;
    end
    if (metaReset) begin
      s2_tag_hit_1 <= 1'h0;
    end else if (s1_valid) begin
      s2_tag_hit_1 <= s1_tag_hit_1;
    end
    if (metaReset) begin
      s2_tag_hit_2 <= 1'h0;
    end else if (s1_valid) begin
      s2_tag_hit_2 <= s1_tag_hit_2;
    end
    if (metaReset) begin
      s2_tag_hit_3 <= 1'h0;
    end else if (s1_valid) begin
      s2_tag_hit_3 <= s1_tag_hit_3;
    end
    if (metaReset) begin
      s2_dout_0 <= 32'h0;
    end else if (s1_valid) begin
      if (io_s1_paddr[2]) begin
        s2_dout_0 <= data_arrays_1_0__T_300_data;
      end else begin
        s2_dout_0 <= _GEN_54;
      end
    end
    if (metaReset) begin
      s2_dout_1 <= 32'h0;
    end else if (s1_valid) begin
      if (io_s1_paddr[2]) begin
        s2_dout_1 <= data_arrays_1_1__T_300_data;
      end else begin
        s2_dout_1 <= _GEN_55;
      end
    end
    if (metaReset) begin
      s2_dout_2 <= 32'h0;
    end else if (s1_valid) begin
      if (io_s1_paddr[2]) begin
        s2_dout_2 <= data_arrays_1_2__T_300_data;
      end else begin
        s2_dout_2 <= _GEN_56;
      end
    end
    if (metaReset) begin
      s2_dout_3 <= 32'h0;
    end else if (s1_valid) begin
      if (io_s1_paddr[2]) begin
        s2_dout_3 <= data_arrays_1_3__T_300_data;
      end else begin
        s2_dout_3 <= _GEN_57;
      end
    end
    if (metaReset) begin
      s2_tl_error <= 1'h0;
    end else if (s1_valid) begin
      s2_tl_error <= _T_329;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_226) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ICache.scala:264 assert(!(s1_valid || s1_slaveValid) || PopCount(s1_tag_hit zip s1_tag_disparity map { case (h, d) => h && !d }) <= 1)\n"); // @[ICache.scala 264:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_226) begin
          $fatal; // @[ICache.scala 264:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    ICache_state <= ICache_xor0;
    if (!(ICache_cov_read_data)) begin
      ICache_covSum <= ICache_covSum + 1'h1;
    end
    if (metaReset) begin
      ICache_metaAssert <= 1'h0;
    end else begin
      ICache_metaAssert <= ICache_metaAssert | ICache_or0;
    end
  end
  always @(posedge clock) begin
    if(ICache_cov_write_en & ICache_cov_write_mask) begin
      ICache_cov[ICache_cov_write_addr] <= ICache_cov_write_data; // @[Coverage map for ICache]
    end
  end
endmodule
module ShiftQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_btb_taken,
  input         io_enq_bits_btb_bridx,
  input  [4:0]  io_enq_bits_btb_entry,
  input  [7:0]  io_enq_bits_btb_bht_history,
  input  [39:0] io_enq_bits_pc,
  input  [31:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_mask,
  input         io_enq_bits_xcpt_pf_inst,
  input         io_enq_bits_xcpt_ae_inst,
  input         io_enq_bits_replay,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_btb_taken,
  output        io_deq_bits_btb_bridx,
  output [4:0]  io_deq_bits_btb_entry,
  output [7:0]  io_deq_bits_btb_bht_history,
  output [39:0] io_deq_bits_pc,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_xcpt_pf_inst,
  output        io_deq_bits_xcpt_ae_inst,
  output        io_deq_bits_replay,
  output [4:0]  io_mask,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  _T_1_0; // @[ShiftQueue.scala 21:30]
  reg [31:0] _RAND_0;
  reg  _T_1_1; // @[ShiftQueue.scala 21:30]
  reg [31:0] _RAND_1;
  reg  _T_1_2; // @[ShiftQueue.scala 21:30]
  reg [31:0] _RAND_2;
  reg  _T_1_3; // @[ShiftQueue.scala 21:30]
  reg [31:0] _RAND_3;
  reg  _T_1_4; // @[ShiftQueue.scala 21:30]
  reg [31:0] _RAND_4;
  reg  _T_2_0_btb_taken; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_5;
  reg  _T_2_0_btb_bridx; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_6;
  reg [4:0] _T_2_0_btb_entry; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_7;
  reg [7:0] _T_2_0_btb_bht_history; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_8;
  reg [39:0] _T_2_0_pc; // @[ShiftQueue.scala 22:25]
  reg [63:0] _RAND_9;
  reg [31:0] _T_2_0_data; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_10;
  reg  _T_2_0_xcpt_pf_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_11;
  reg  _T_2_0_xcpt_ae_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_12;
  reg  _T_2_0_replay; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_13;
  reg  _T_2_1_btb_taken; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_14;
  reg  _T_2_1_btb_bridx; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_15;
  reg [4:0] _T_2_1_btb_entry; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_16;
  reg [7:0] _T_2_1_btb_bht_history; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_17;
  reg [39:0] _T_2_1_pc; // @[ShiftQueue.scala 22:25]
  reg [63:0] _RAND_18;
  reg [31:0] _T_2_1_data; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_19;
  reg  _T_2_1_xcpt_pf_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_20;
  reg  _T_2_1_xcpt_ae_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_21;
  reg  _T_2_1_replay; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_22;
  reg  _T_2_2_btb_taken; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_23;
  reg  _T_2_2_btb_bridx; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_24;
  reg [4:0] _T_2_2_btb_entry; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_25;
  reg [7:0] _T_2_2_btb_bht_history; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_26;
  reg [39:0] _T_2_2_pc; // @[ShiftQueue.scala 22:25]
  reg [63:0] _RAND_27;
  reg [31:0] _T_2_2_data; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_28;
  reg  _T_2_2_xcpt_pf_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_29;
  reg  _T_2_2_xcpt_ae_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_30;
  reg  _T_2_2_replay; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_31;
  reg  _T_2_3_btb_taken; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_32;
  reg  _T_2_3_btb_bridx; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_33;
  reg [4:0] _T_2_3_btb_entry; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_34;
  reg [7:0] _T_2_3_btb_bht_history; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_35;
  reg [39:0] _T_2_3_pc; // @[ShiftQueue.scala 22:25]
  reg [63:0] _RAND_36;
  reg [31:0] _T_2_3_data; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_37;
  reg  _T_2_3_xcpt_pf_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_38;
  reg  _T_2_3_xcpt_ae_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_39;
  reg  _T_2_3_replay; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_40;
  reg  _T_2_4_btb_taken; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_41;
  reg  _T_2_4_btb_bridx; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_42;
  reg [4:0] _T_2_4_btb_entry; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_43;
  reg [7:0] _T_2_4_btb_bht_history; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_44;
  reg [39:0] _T_2_4_pc; // @[ShiftQueue.scala 22:25]
  reg [63:0] _RAND_45;
  reg [31:0] _T_2_4_data; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_46;
  reg  _T_2_4_xcpt_pf_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_47;
  reg  _T_2_4_xcpt_ae_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_48;
  reg  _T_2_4_replay; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_49;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[ShiftQueue.scala 30:45]
  wire  _T_7; // @[ShiftQueue.scala 30:28]
  wire  _T_11; // @[ShiftQueue.scala 31:45]
  wire  _T_12; // @[ShiftQueue.scala 29:10]
  wire  _T_19; // @[ShiftQueue.scala 37:45]
  wire  _T_24; // @[ShiftQueue.scala 30:45]
  wire  _T_25; // @[ShiftQueue.scala 30:28]
  wire  _T_29; // @[ShiftQueue.scala 31:45]
  wire  _T_30; // @[ShiftQueue.scala 29:10]
  wire  _T_37; // @[ShiftQueue.scala 37:45]
  wire  _T_42; // @[ShiftQueue.scala 30:45]
  wire  _T_43; // @[ShiftQueue.scala 30:28]
  wire  _T_47; // @[ShiftQueue.scala 31:45]
  wire  _T_48; // @[ShiftQueue.scala 29:10]
  wire  _T_55; // @[ShiftQueue.scala 37:45]
  wire  _T_60; // @[ShiftQueue.scala 30:45]
  wire  _T_61; // @[ShiftQueue.scala 30:28]
  wire  _T_65; // @[ShiftQueue.scala 31:45]
  wire  _T_66; // @[ShiftQueue.scala 29:10]
  wire  _T_73; // @[ShiftQueue.scala 37:45]
  wire  _T_77; // @[ShiftQueue.scala 30:45]
  wire  _T_82; // @[ShiftQueue.scala 31:45]
  wire  _T_83; // @[ShiftQueue.scala 29:10]
  wire  _T_90; // @[ShiftQueue.scala 37:45]
  wire [1:0] _T_94; // @[ShiftQueue.scala 53:20]
  wire [2:0] _T_96; // @[ShiftQueue.scala 53:20]
  reg  ShiftQueue_state; // @[Register tracking ShiftQueue state]
  reg [31:0] _RAND_50;
  reg  ShiftQueue_cov [0:1]; // @[Coverage map for ShiftQueue]
  reg [31:0] _RAND_51;
  wire  ShiftQueue_cov_read_data; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_read_addr; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_write_data; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_write_addr; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_write_mask; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_write_en; // @[Coverage map for ShiftQueue]
  reg [29:0] ShiftQueue_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_52;
  wire  _T_1_4_shl;
  wire  _T_1_4_pad;
  wire  _T_1_1_shl;
  wire  _T_1_1_pad;
  wire  _T_1_2_shl;
  wire  _T_1_2_pad;
  wire  _T_1_0_shl;
  wire  _T_1_0_pad;
  wire  _T_1_3_shl;
  wire  _T_1_3_pad;
  wire  ShiftQueue_xor1;
  wire  ShiftQueue_xor6;
  wire  ShiftQueue_xor2;
  wire  ShiftQueue_xor0;
  assign _T_4 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = _T_4 & _T_1_0; // @[ShiftQueue.scala 30:45]
  assign _T_7 = _T_1_1 | _T_6; // @[ShiftQueue.scala 30:28]
  assign _T_11 = _T_4 & ~_T_1_0; // @[ShiftQueue.scala 31:45]
  assign _T_12 = io_deq_ready ? _T_7 : _T_11; // @[ShiftQueue.scala 29:10]
  assign _T_19 = _T_4 | _T_1_0; // @[ShiftQueue.scala 37:45]
  assign _T_24 = _T_4 & _T_1_1; // @[ShiftQueue.scala 30:45]
  assign _T_25 = _T_1_2 | _T_24; // @[ShiftQueue.scala 30:28]
  assign _T_29 = _T_6 & ~_T_1_1; // @[ShiftQueue.scala 31:45]
  assign _T_30 = io_deq_ready ? _T_25 : _T_29; // @[ShiftQueue.scala 29:10]
  assign _T_37 = _T_6 | _T_1_1; // @[ShiftQueue.scala 37:45]
  assign _T_42 = _T_4 & _T_1_2; // @[ShiftQueue.scala 30:45]
  assign _T_43 = _T_1_3 | _T_42; // @[ShiftQueue.scala 30:28]
  assign _T_47 = _T_24 & ~_T_1_2; // @[ShiftQueue.scala 31:45]
  assign _T_48 = io_deq_ready ? _T_43 : _T_47; // @[ShiftQueue.scala 29:10]
  assign _T_55 = _T_24 | _T_1_2; // @[ShiftQueue.scala 37:45]
  assign _T_60 = _T_4 & _T_1_3; // @[ShiftQueue.scala 30:45]
  assign _T_61 = _T_1_4 | _T_60; // @[ShiftQueue.scala 30:28]
  assign _T_65 = _T_42 & ~_T_1_3; // @[ShiftQueue.scala 31:45]
  assign _T_66 = io_deq_ready ? _T_61 : _T_65; // @[ShiftQueue.scala 29:10]
  assign _T_73 = _T_42 | _T_1_3; // @[ShiftQueue.scala 37:45]
  assign _T_77 = _T_4 & _T_1_4; // @[ShiftQueue.scala 30:45]
  assign _T_82 = _T_60 & ~_T_1_4; // @[ShiftQueue.scala 31:45]
  assign _T_83 = io_deq_ready ? _T_77 : _T_82; // @[ShiftQueue.scala 29:10]
  assign _T_90 = _T_60 | _T_1_4; // @[ShiftQueue.scala 37:45]
  assign _T_94 = {_T_1_1,_T_1_0}; // @[ShiftQueue.scala 53:20]
  assign _T_96 = {_T_1_4,_T_1_3,_T_1_2}; // @[ShiftQueue.scala 53:20]
  assign io_enq_ready = ~_T_1_4; // @[ShiftQueue.scala 40:16]
  assign io_deq_valid = io_enq_valid | _T_1_0; // @[ShiftQueue.scala 41:16 ShiftQueue.scala 45:40]
  assign io_deq_bits_btb_taken = _T_1_0 ? _T_2_0_btb_taken : io_enq_bits_btb_taken; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_btb_bridx = _T_1_0 ? _T_2_0_btb_bridx : io_enq_bits_btb_bridx; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_btb_entry = _T_1_0 ? _T_2_0_btb_entry : io_enq_bits_btb_entry; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_btb_bht_history = _T_1_0 ? _T_2_0_btb_bht_history : io_enq_bits_btb_bht_history; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_pc = _T_1_0 ? _T_2_0_pc : io_enq_bits_pc; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_data = _T_1_0 ? _T_2_0_data : io_enq_bits_data; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_xcpt_pf_inst = _T_1_0 ? _T_2_0_xcpt_pf_inst : io_enq_bits_xcpt_pf_inst; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_xcpt_ae_inst = _T_1_0 ? _T_2_0_xcpt_ae_inst : io_enq_bits_xcpt_ae_inst; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_replay = _T_1_0 ? _T_2_0_replay : io_enq_bits_replay; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_mask = {_T_96,_T_94}; // @[ShiftQueue.scala 53:11]
  assign ShiftQueue_cov_read_addr = ShiftQueue_state;
  assign ShiftQueue_cov_read_data = ShiftQueue_cov[ShiftQueue_cov_read_addr]; // @[Coverage map for ShiftQueue]
  assign ShiftQueue_cov_write_data = 1'h1;
  assign ShiftQueue_cov_write_addr = ShiftQueue_state;
  assign ShiftQueue_cov_write_mask = 1'h1;
  assign ShiftQueue_cov_write_en = 1'h1;
  assign _T_1_4_shl = _T_1_4;
  assign _T_1_4_pad = _T_1_4_shl;
  assign _T_1_1_shl = _T_1_1;
  assign _T_1_1_pad = _T_1_1_shl;
  assign _T_1_2_shl = _T_1_2;
  assign _T_1_2_pad = _T_1_2_shl;
  assign _T_1_0_shl = _T_1_0;
  assign _T_1_0_pad = _T_1_0_shl;
  assign _T_1_3_shl = _T_1_3;
  assign _T_1_3_pad = _T_1_3_shl;
  assign ShiftQueue_xor1 = _T_1_4_pad ^ _T_1_1_pad;
  assign ShiftQueue_xor6 = _T_1_0_pad ^ _T_1_3_pad;
  assign ShiftQueue_xor2 = _T_1_2_pad ^ ShiftQueue_xor6;
  assign ShiftQueue_xor0 = ShiftQueue_xor1 ^ ShiftQueue_xor2;
  assign io_covSum = ShiftQueue_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2_0_btb_taken = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2_0_btb_bridx = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2_0_btb_entry = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2_0_btb_bht_history = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  _T_2_0_pc = _RAND_9[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2_0_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2_0_xcpt_pf_inst = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2_0_xcpt_ae_inst = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2_0_replay = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_2_1_btb_taken = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2_1_btb_bridx = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_2_1_btb_entry = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_2_1_btb_bht_history = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  _T_2_1_pc = _RAND_18[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_2_1_data = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_2_1_xcpt_pf_inst = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_2_1_xcpt_ae_inst = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_2_1_replay = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_2_2_btb_taken = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_2_2_btb_bridx = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_2_2_btb_entry = _RAND_25[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_2_2_btb_bht_history = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  _T_2_2_pc = _RAND_27[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_2_2_data = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_2_2_xcpt_pf_inst = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_2_2_xcpt_ae_inst = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_2_2_replay = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_2_3_btb_taken = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_2_3_btb_bridx = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_2_3_btb_entry = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_2_3_btb_bht_history = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{`RANDOM}};
  _T_2_3_pc = _RAND_36[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_2_3_data = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_2_3_xcpt_pf_inst = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_2_3_xcpt_ae_inst = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_2_3_replay = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_2_4_btb_taken = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_2_4_btb_bridx = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_2_4_btb_entry = _RAND_43[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_2_4_btb_bht_history = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {2{`RANDOM}};
  _T_2_4_pc = _RAND_45[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_2_4_data = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_2_4_xcpt_pf_inst = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_2_4_xcpt_ae_inst = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_2_4_replay = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  ShiftQueue_state = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ShiftQueue_cov[initvar] = _RAND_51[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  ShiftQueue_covSum = _RAND_52[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_1_0 <= 1'h0;
    end else if (reset) begin
      _T_1_0 <= 1'h0;
    end else if (io_deq_ready) begin
      _T_1_0 <= _T_7;
    end else begin
      _T_1_0 <= _T_19;
    end
    if (metaReset) begin
      _T_1_1 <= 1'h0;
    end else if (reset) begin
      _T_1_1 <= 1'h0;
    end else if (io_deq_ready) begin
      _T_1_1 <= _T_25;
    end else begin
      _T_1_1 <= _T_37;
    end
    if (metaReset) begin
      _T_1_2 <= 1'h0;
    end else if (reset) begin
      _T_1_2 <= 1'h0;
    end else if (io_deq_ready) begin
      _T_1_2 <= _T_43;
    end else begin
      _T_1_2 <= _T_55;
    end
    if (metaReset) begin
      _T_1_3 <= 1'h0;
    end else if (reset) begin
      _T_1_3 <= 1'h0;
    end else if (io_deq_ready) begin
      _T_1_3 <= _T_61;
    end else begin
      _T_1_3 <= _T_73;
    end
    if (metaReset) begin
      _T_1_4 <= 1'h0;
    end else if (reset) begin
      _T_1_4 <= 1'h0;
    end else if (io_deq_ready) begin
      _T_1_4 <= _T_77;
    end else begin
      _T_1_4 <= _T_90;
    end
    if (metaReset) begin
      _T_2_0_btb_taken <= 1'h0;
    end else if (_T_12) begin
      if (_T_1_1) begin
        _T_2_0_btb_taken <= _T_2_1_btb_taken;
      end else begin
        _T_2_0_btb_taken <= io_enq_bits_btb_taken;
      end
    end
    if (metaReset) begin
      _T_2_0_btb_bridx <= 1'h0;
    end else if (_T_12) begin
      if (_T_1_1) begin
        _T_2_0_btb_bridx <= _T_2_1_btb_bridx;
      end else begin
        _T_2_0_btb_bridx <= io_enq_bits_btb_bridx;
      end
    end
    if (metaReset) begin
      _T_2_0_btb_entry <= 5'h0;
    end else if (_T_12) begin
      if (_T_1_1) begin
        _T_2_0_btb_entry <= _T_2_1_btb_entry;
      end else begin
        _T_2_0_btb_entry <= io_enq_bits_btb_entry;
      end
    end
    if (metaReset) begin
      _T_2_0_btb_bht_history <= 8'h0;
    end else if (_T_12) begin
      if (_T_1_1) begin
        _T_2_0_btb_bht_history <= _T_2_1_btb_bht_history;
      end else begin
        _T_2_0_btb_bht_history <= io_enq_bits_btb_bht_history;
      end
    end
    if (metaReset) begin
      _T_2_0_pc <= 40'h0;
    end else if (_T_12) begin
      if (_T_1_1) begin
        _T_2_0_pc <= _T_2_1_pc;
      end else begin
        _T_2_0_pc <= io_enq_bits_pc;
      end
    end
    if (metaReset) begin
      _T_2_0_data <= 32'h0;
    end else if (_T_12) begin
      if (_T_1_1) begin
        _T_2_0_data <= _T_2_1_data;
      end else begin
        _T_2_0_data <= io_enq_bits_data;
      end
    end
    if (metaReset) begin
      _T_2_0_xcpt_pf_inst <= 1'h0;
    end else if (_T_12) begin
      if (_T_1_1) begin
        _T_2_0_xcpt_pf_inst <= _T_2_1_xcpt_pf_inst;
      end else begin
        _T_2_0_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      _T_2_0_xcpt_ae_inst <= 1'h0;
    end else if (_T_12) begin
      if (_T_1_1) begin
        _T_2_0_xcpt_ae_inst <= _T_2_1_xcpt_ae_inst;
      end else begin
        _T_2_0_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      _T_2_0_replay <= 1'h0;
    end else if (_T_12) begin
      if (_T_1_1) begin
        _T_2_0_replay <= _T_2_1_replay;
      end else begin
        _T_2_0_replay <= io_enq_bits_replay;
      end
    end
    if (metaReset) begin
      _T_2_1_btb_taken <= 1'h0;
    end else if (_T_30) begin
      if (_T_1_2) begin
        _T_2_1_btb_taken <= _T_2_2_btb_taken;
      end else begin
        _T_2_1_btb_taken <= io_enq_bits_btb_taken;
      end
    end
    if (metaReset) begin
      _T_2_1_btb_bridx <= 1'h0;
    end else if (_T_30) begin
      if (_T_1_2) begin
        _T_2_1_btb_bridx <= _T_2_2_btb_bridx;
      end else begin
        _T_2_1_btb_bridx <= io_enq_bits_btb_bridx;
      end
    end
    if (metaReset) begin
      _T_2_1_btb_entry <= 5'h0;
    end else if (_T_30) begin
      if (_T_1_2) begin
        _T_2_1_btb_entry <= _T_2_2_btb_entry;
      end else begin
        _T_2_1_btb_entry <= io_enq_bits_btb_entry;
      end
    end
    if (metaReset) begin
      _T_2_1_btb_bht_history <= 8'h0;
    end else if (_T_30) begin
      if (_T_1_2) begin
        _T_2_1_btb_bht_history <= _T_2_2_btb_bht_history;
      end else begin
        _T_2_1_btb_bht_history <= io_enq_bits_btb_bht_history;
      end
    end
    if (metaReset) begin
      _T_2_1_pc <= 40'h0;
    end else if (_T_30) begin
      if (_T_1_2) begin
        _T_2_1_pc <= _T_2_2_pc;
      end else begin
        _T_2_1_pc <= io_enq_bits_pc;
      end
    end
    if (metaReset) begin
      _T_2_1_data <= 32'h0;
    end else if (_T_30) begin
      if (_T_1_2) begin
        _T_2_1_data <= _T_2_2_data;
      end else begin
        _T_2_1_data <= io_enq_bits_data;
      end
    end
    if (metaReset) begin
      _T_2_1_xcpt_pf_inst <= 1'h0;
    end else if (_T_30) begin
      if (_T_1_2) begin
        _T_2_1_xcpt_pf_inst <= _T_2_2_xcpt_pf_inst;
      end else begin
        _T_2_1_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      _T_2_1_xcpt_ae_inst <= 1'h0;
    end else if (_T_30) begin
      if (_T_1_2) begin
        _T_2_1_xcpt_ae_inst <= _T_2_2_xcpt_ae_inst;
      end else begin
        _T_2_1_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      _T_2_1_replay <= 1'h0;
    end else if (_T_30) begin
      if (_T_1_2) begin
        _T_2_1_replay <= _T_2_2_replay;
      end else begin
        _T_2_1_replay <= io_enq_bits_replay;
      end
    end
    if (metaReset) begin
      _T_2_2_btb_taken <= 1'h0;
    end else if (_T_48) begin
      if (_T_1_3) begin
        _T_2_2_btb_taken <= _T_2_3_btb_taken;
      end else begin
        _T_2_2_btb_taken <= io_enq_bits_btb_taken;
      end
    end
    if (metaReset) begin
      _T_2_2_btb_bridx <= 1'h0;
    end else if (_T_48) begin
      if (_T_1_3) begin
        _T_2_2_btb_bridx <= _T_2_3_btb_bridx;
      end else begin
        _T_2_2_btb_bridx <= io_enq_bits_btb_bridx;
      end
    end
    if (metaReset) begin
      _T_2_2_btb_entry <= 5'h0;
    end else if (_T_48) begin
      if (_T_1_3) begin
        _T_2_2_btb_entry <= _T_2_3_btb_entry;
      end else begin
        _T_2_2_btb_entry <= io_enq_bits_btb_entry;
      end
    end
    if (metaReset) begin
      _T_2_2_btb_bht_history <= 8'h0;
    end else if (_T_48) begin
      if (_T_1_3) begin
        _T_2_2_btb_bht_history <= _T_2_3_btb_bht_history;
      end else begin
        _T_2_2_btb_bht_history <= io_enq_bits_btb_bht_history;
      end
    end
    if (metaReset) begin
      _T_2_2_pc <= 40'h0;
    end else if (_T_48) begin
      if (_T_1_3) begin
        _T_2_2_pc <= _T_2_3_pc;
      end else begin
        _T_2_2_pc <= io_enq_bits_pc;
      end
    end
    if (metaReset) begin
      _T_2_2_data <= 32'h0;
    end else if (_T_48) begin
      if (_T_1_3) begin
        _T_2_2_data <= _T_2_3_data;
      end else begin
        _T_2_2_data <= io_enq_bits_data;
      end
    end
    if (metaReset) begin
      _T_2_2_xcpt_pf_inst <= 1'h0;
    end else if (_T_48) begin
      if (_T_1_3) begin
        _T_2_2_xcpt_pf_inst <= _T_2_3_xcpt_pf_inst;
      end else begin
        _T_2_2_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      _T_2_2_xcpt_ae_inst <= 1'h0;
    end else if (_T_48) begin
      if (_T_1_3) begin
        _T_2_2_xcpt_ae_inst <= _T_2_3_xcpt_ae_inst;
      end else begin
        _T_2_2_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      _T_2_2_replay <= 1'h0;
    end else if (_T_48) begin
      if (_T_1_3) begin
        _T_2_2_replay <= _T_2_3_replay;
      end else begin
        _T_2_2_replay <= io_enq_bits_replay;
      end
    end
    if (metaReset) begin
      _T_2_3_btb_taken <= 1'h0;
    end else if (_T_66) begin
      if (_T_1_4) begin
        _T_2_3_btb_taken <= _T_2_4_btb_taken;
      end else begin
        _T_2_3_btb_taken <= io_enq_bits_btb_taken;
      end
    end
    if (metaReset) begin
      _T_2_3_btb_bridx <= 1'h0;
    end else if (_T_66) begin
      if (_T_1_4) begin
        _T_2_3_btb_bridx <= _T_2_4_btb_bridx;
      end else begin
        _T_2_3_btb_bridx <= io_enq_bits_btb_bridx;
      end
    end
    if (metaReset) begin
      _T_2_3_btb_entry <= 5'h0;
    end else if (_T_66) begin
      if (_T_1_4) begin
        _T_2_3_btb_entry <= _T_2_4_btb_entry;
      end else begin
        _T_2_3_btb_entry <= io_enq_bits_btb_entry;
      end
    end
    if (metaReset) begin
      _T_2_3_btb_bht_history <= 8'h0;
    end else if (_T_66) begin
      if (_T_1_4) begin
        _T_2_3_btb_bht_history <= _T_2_4_btb_bht_history;
      end else begin
        _T_2_3_btb_bht_history <= io_enq_bits_btb_bht_history;
      end
    end
    if (metaReset) begin
      _T_2_3_pc <= 40'h0;
    end else if (_T_66) begin
      if (_T_1_4) begin
        _T_2_3_pc <= _T_2_4_pc;
      end else begin
        _T_2_3_pc <= io_enq_bits_pc;
      end
    end
    if (metaReset) begin
      _T_2_3_data <= 32'h0;
    end else if (_T_66) begin
      if (_T_1_4) begin
        _T_2_3_data <= _T_2_4_data;
      end else begin
        _T_2_3_data <= io_enq_bits_data;
      end
    end
    if (metaReset) begin
      _T_2_3_xcpt_pf_inst <= 1'h0;
    end else if (_T_66) begin
      if (_T_1_4) begin
        _T_2_3_xcpt_pf_inst <= _T_2_4_xcpt_pf_inst;
      end else begin
        _T_2_3_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      _T_2_3_xcpt_ae_inst <= 1'h0;
    end else if (_T_66) begin
      if (_T_1_4) begin
        _T_2_3_xcpt_ae_inst <= _T_2_4_xcpt_ae_inst;
      end else begin
        _T_2_3_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      _T_2_3_replay <= 1'h0;
    end else if (_T_66) begin
      if (_T_1_4) begin
        _T_2_3_replay <= _T_2_4_replay;
      end else begin
        _T_2_3_replay <= io_enq_bits_replay;
      end
    end
    if (metaReset) begin
      _T_2_4_btb_taken <= 1'h0;
    end else if (_T_83) begin
      _T_2_4_btb_taken <= io_enq_bits_btb_taken;
    end
    if (metaReset) begin
      _T_2_4_btb_bridx <= 1'h0;
    end else if (_T_83) begin
      _T_2_4_btb_bridx <= io_enq_bits_btb_bridx;
    end
    if (metaReset) begin
      _T_2_4_btb_entry <= 5'h0;
    end else if (_T_83) begin
      _T_2_4_btb_entry <= io_enq_bits_btb_entry;
    end
    if (metaReset) begin
      _T_2_4_btb_bht_history <= 8'h0;
    end else if (_T_83) begin
      _T_2_4_btb_bht_history <= io_enq_bits_btb_bht_history;
    end
    if (metaReset) begin
      _T_2_4_pc <= 40'h0;
    end else if (_T_83) begin
      _T_2_4_pc <= io_enq_bits_pc;
    end
    if (metaReset) begin
      _T_2_4_data <= 32'h0;
    end else if (_T_83) begin
      _T_2_4_data <= io_enq_bits_data;
    end
    if (metaReset) begin
      _T_2_4_xcpt_pf_inst <= 1'h0;
    end else if (_T_83) begin
      _T_2_4_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
    end
    if (metaReset) begin
      _T_2_4_xcpt_ae_inst <= 1'h0;
    end else if (_T_83) begin
      _T_2_4_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
    end
    if (metaReset) begin
      _T_2_4_replay <= 1'h0;
    end else if (_T_83) begin
      _T_2_4_replay <= io_enq_bits_replay;
    end
    ShiftQueue_state <= ShiftQueue_xor0;
    if (!(ShiftQueue_cov_read_data)) begin
      ShiftQueue_covSum <= ShiftQueue_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(ShiftQueue_cov_write_en & ShiftQueue_cov_write_mask) begin
      ShiftQueue_cov[ShiftQueue_cov_write_addr] <= ShiftQueue_cov_write_data; // @[Coverage map for ShiftQueue]
    end
  end
endmodule
module TLB_1(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [39:0] io_req_bits_vaddr,
  output        io_resp_miss,
  output [31:0] io_resp_paddr,
  output        io_resp_pf_inst,
  output        io_resp_ae_inst,
  output        io_resp_cacheable,
  input         io_sfence_valid,
  input         io_sfence_bits_rs1,
  input         io_sfence_bits_rs2,
  input  [38:0] io_sfence_bits_addr,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output        io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input         io_ptw_status_debug,
  input  [1:0]  io_ptw_status_prv,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input         io_kill,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [19:0] OptimizationBarrier_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_metaAssert; // @[package.scala 236:25]
  wire [1:0] pmp_io_prv; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_0_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_0_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_1_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_1_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_2_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_2_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_3_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_3_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_4_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_4_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_5_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_5_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_6_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_6_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_7_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_7_mask; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_addr; // @[TLB.scala 190:19]
  wire  pmp_io_r; // @[TLB.scala 190:19]
  wire  pmp_io_w; // @[TLB.scala 190:19]
  wire  pmp_io_x; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_covSum; // @[TLB.scala 190:19]
  wire  pmp_metaAssert; // @[TLB.scala 190:19]
  wire [19:0] OptimizationBarrier_1_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_1_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_1_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_1_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_2_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_2_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_2_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_2_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_3_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_3_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_3_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_3_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_4_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_4_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_4_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_4_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_5_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_5_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_5_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_5_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_6_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_6_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_6_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_6_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_7_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_7_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_7_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_7_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_8_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_8_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_8_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_8_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_9_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_9_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_9_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_9_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_10_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_10_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_10_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_10_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_11_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_11_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_11_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_11_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_12_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_12_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_12_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_12_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_13_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_13_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_13_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_13_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_14_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_14_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_14_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_14_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_15_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_15_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_15_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_15_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_16_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_16_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_16_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_16_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_17_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_17_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_17_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_17_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_18_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_18_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_18_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_18_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_19_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_19_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_19_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_19_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_20_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_20_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_20_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_20_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_21_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_21_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_21_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_21_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_22_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_22_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_22_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_22_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_23_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_23_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_23_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_23_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_24_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_24_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_24_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_24_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_25_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_25_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_25_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_25_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_26_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_26_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_26_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_26_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_27_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_27_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_27_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_27_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_28_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_28_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_28_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_28_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_29_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_29_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_29_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_29_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_30_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_30_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_30_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_30_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_31_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_31_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_31_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_31_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_32_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_32_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_32_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_32_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_33_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_33_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_33_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_33_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_34_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_34_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_34_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_34_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_35_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_35_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_35_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_35_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_36_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_36_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_36_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_36_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_37_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_37_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_37_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_37_metaAssert; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_38_io_x_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_x_c; // @[package.scala 236:25]
  wire [19:0] OptimizationBarrier_38_io_y_ppn; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_u; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_ae; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_sw; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_sx; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_sr; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_pw; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_px; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_pr; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_ppp; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_pal; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_paa; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_eff; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_io_y_c; // @[package.scala 236:25]
  wire [29:0] OptimizationBarrier_38_io_covSum; // @[package.scala 236:25]
  wire  OptimizationBarrier_38_metaAssert; // @[package.scala 236:25]
  reg [26:0] sectored_entries_0_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_0;
  reg [34:0] sectored_entries_0_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_1;
  reg [34:0] sectored_entries_0_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_2;
  reg [34:0] sectored_entries_0_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_3;
  reg [34:0] sectored_entries_0_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_4;
  reg  sectored_entries_0_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_5;
  reg  sectored_entries_0_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_6;
  reg  sectored_entries_0_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_7;
  reg  sectored_entries_0_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_8;
  reg [26:0] sectored_entries_1_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_9;
  reg [34:0] sectored_entries_1_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_10;
  reg [34:0] sectored_entries_1_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_11;
  reg [34:0] sectored_entries_1_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_12;
  reg [34:0] sectored_entries_1_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_13;
  reg  sectored_entries_1_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_14;
  reg  sectored_entries_1_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_15;
  reg  sectored_entries_1_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_16;
  reg  sectored_entries_1_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_17;
  reg [26:0] sectored_entries_2_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_18;
  reg [34:0] sectored_entries_2_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_19;
  reg [34:0] sectored_entries_2_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_20;
  reg [34:0] sectored_entries_2_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_21;
  reg [34:0] sectored_entries_2_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_22;
  reg  sectored_entries_2_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_23;
  reg  sectored_entries_2_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_24;
  reg  sectored_entries_2_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_25;
  reg  sectored_entries_2_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_26;
  reg [26:0] sectored_entries_3_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_27;
  reg [34:0] sectored_entries_3_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_28;
  reg [34:0] sectored_entries_3_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_29;
  reg [34:0] sectored_entries_3_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_30;
  reg [34:0] sectored_entries_3_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_31;
  reg  sectored_entries_3_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_32;
  reg  sectored_entries_3_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_33;
  reg  sectored_entries_3_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_34;
  reg  sectored_entries_3_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_35;
  reg [26:0] sectored_entries_4_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_36;
  reg [34:0] sectored_entries_4_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_37;
  reg [34:0] sectored_entries_4_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_38;
  reg [34:0] sectored_entries_4_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_39;
  reg [34:0] sectored_entries_4_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_40;
  reg  sectored_entries_4_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_41;
  reg  sectored_entries_4_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_42;
  reg  sectored_entries_4_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_43;
  reg  sectored_entries_4_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_44;
  reg [26:0] sectored_entries_5_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_45;
  reg [34:0] sectored_entries_5_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_46;
  reg [34:0] sectored_entries_5_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_47;
  reg [34:0] sectored_entries_5_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_48;
  reg [34:0] sectored_entries_5_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_49;
  reg  sectored_entries_5_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_50;
  reg  sectored_entries_5_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_51;
  reg  sectored_entries_5_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_52;
  reg  sectored_entries_5_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_53;
  reg [26:0] sectored_entries_6_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_54;
  reg [34:0] sectored_entries_6_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_55;
  reg [34:0] sectored_entries_6_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_56;
  reg [34:0] sectored_entries_6_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_57;
  reg [34:0] sectored_entries_6_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_58;
  reg  sectored_entries_6_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_59;
  reg  sectored_entries_6_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_60;
  reg  sectored_entries_6_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_61;
  reg  sectored_entries_6_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_62;
  reg [26:0] sectored_entries_7_tag; // @[TLB.scala 162:29]
  reg [31:0] _RAND_63;
  reg [34:0] sectored_entries_7_data_0; // @[TLB.scala 162:29]
  reg [63:0] _RAND_64;
  reg [34:0] sectored_entries_7_data_1; // @[TLB.scala 162:29]
  reg [63:0] _RAND_65;
  reg [34:0] sectored_entries_7_data_2; // @[TLB.scala 162:29]
  reg [63:0] _RAND_66;
  reg [34:0] sectored_entries_7_data_3; // @[TLB.scala 162:29]
  reg [63:0] _RAND_67;
  reg  sectored_entries_7_valid_0; // @[TLB.scala 162:29]
  reg [31:0] _RAND_68;
  reg  sectored_entries_7_valid_1; // @[TLB.scala 162:29]
  reg [31:0] _RAND_69;
  reg  sectored_entries_7_valid_2; // @[TLB.scala 162:29]
  reg [31:0] _RAND_70;
  reg  sectored_entries_7_valid_3; // @[TLB.scala 162:29]
  reg [31:0] _RAND_71;
  reg [1:0] superpage_entries_0_level; // @[TLB.scala 163:30]
  reg [31:0] _RAND_72;
  reg [26:0] superpage_entries_0_tag; // @[TLB.scala 163:30]
  reg [31:0] _RAND_73;
  reg [34:0] superpage_entries_0_data_0; // @[TLB.scala 163:30]
  reg [63:0] _RAND_74;
  reg  superpage_entries_0_valid_0; // @[TLB.scala 163:30]
  reg [31:0] _RAND_75;
  reg [1:0] superpage_entries_1_level; // @[TLB.scala 163:30]
  reg [31:0] _RAND_76;
  reg [26:0] superpage_entries_1_tag; // @[TLB.scala 163:30]
  reg [31:0] _RAND_77;
  reg [34:0] superpage_entries_1_data_0; // @[TLB.scala 163:30]
  reg [63:0] _RAND_78;
  reg  superpage_entries_1_valid_0; // @[TLB.scala 163:30]
  reg [31:0] _RAND_79;
  reg [1:0] superpage_entries_2_level; // @[TLB.scala 163:30]
  reg [31:0] _RAND_80;
  reg [26:0] superpage_entries_2_tag; // @[TLB.scala 163:30]
  reg [31:0] _RAND_81;
  reg [34:0] superpage_entries_2_data_0; // @[TLB.scala 163:30]
  reg [63:0] _RAND_82;
  reg  superpage_entries_2_valid_0; // @[TLB.scala 163:30]
  reg [31:0] _RAND_83;
  reg [1:0] superpage_entries_3_level; // @[TLB.scala 163:30]
  reg [31:0] _RAND_84;
  reg [26:0] superpage_entries_3_tag; // @[TLB.scala 163:30]
  reg [31:0] _RAND_85;
  reg [34:0] superpage_entries_3_data_0; // @[TLB.scala 163:30]
  reg [63:0] _RAND_86;
  reg  superpage_entries_3_valid_0; // @[TLB.scala 163:30]
  reg [31:0] _RAND_87;
  reg [1:0] special_entry_level; // @[TLB.scala 164:56]
  reg [31:0] _RAND_88;
  reg [26:0] special_entry_tag; // @[TLB.scala 164:56]
  reg [31:0] _RAND_89;
  reg [34:0] special_entry_data_0; // @[TLB.scala 164:56]
  reg [63:0] _RAND_90;
  reg  special_entry_valid_0; // @[TLB.scala 164:56]
  reg [31:0] _RAND_91;
  reg [1:0] state; // @[TLB.scala 169:18]
  reg [31:0] _RAND_92;
  reg [26:0] r_refill_tag; // @[TLB.scala 170:25]
  reg [31:0] _RAND_93;
  reg [1:0] r_superpage_repl_addr; // @[TLB.scala 171:34]
  reg [31:0] _RAND_94;
  reg [2:0] r_sectored_repl_addr; // @[TLB.scala 172:33]
  reg [31:0] _RAND_95;
  reg [2:0] r_sectored_hit_addr; // @[TLB.scala 173:32]
  reg [31:0] _RAND_96;
  reg  r_sectored_hit; // @[TLB.scala 174:27]
  reg [31:0] _RAND_97;
  wire  priv_s; // @[TLB.scala 177:20]
  wire  priv_uses_vm; // @[TLB.scala 178:27]
  wire  vm_enabled; // @[TLB.scala 179:83]
  wire [26:0] vpn; // @[TLB.scala 182:30]
  wire [19:0] refill_ppn; // @[TLB.scala 183:44]
  wire  _T_4; // @[package.scala 15:47]
  wire  _T_5; // @[package.scala 15:47]
  wire  _T_6; // @[package.scala 64:59]
  wire  invalidate_refill; // @[TLB.scala 185:88]
  wire  _T_27; // @[TLB.scala 108:28]
  wire [26:0] _T_29; // @[TLB.scala 109:28]
  wire [26:0] _GEN_983; // @[TLB.scala 109:47]
  wire [26:0] _T_30; // @[TLB.scala 109:47]
  wire  _T_33; // @[TLB.scala 108:28]
  wire [26:0] _T_35; // @[TLB.scala 109:28]
  wire [26:0] _T_36; // @[TLB.scala 109:47]
  wire [19:0] _T_38; // @[Cat.scala 29:58]
  wire [27:0] _T_40; // @[TLB.scala 187:20]
  wire [27:0] mpu_ppn; // @[TLB.scala 186:20]
  wire [39:0] mpu_physaddr; // @[Cat.scala 29:58]
  wire [2:0] _T_44; // @[Cat.scala 29:58]
  wire [2:0] mpu_priv; // @[TLB.scala 189:27]
  wire [39:0] _T_45; // @[Parameters.scala 137:31]
  wire [40:0] _T_46; // @[Parameters.scala 137:49]
  wire [40:0] _T_48; // @[Parameters.scala 137:52]
  wire  _T_49; // @[Parameters.scala 137:67]
  wire [39:0] _T_50; // @[Parameters.scala 137:31]
  wire [40:0] _T_51; // @[Parameters.scala 137:49]
  wire [40:0] _T_53; // @[Parameters.scala 137:52]
  wire  _T_54; // @[Parameters.scala 137:67]
  wire [39:0] _T_55; // @[Parameters.scala 137:31]
  wire [40:0] _T_56; // @[Parameters.scala 137:49]
  wire [40:0] _T_58; // @[Parameters.scala 137:52]
  wire  _T_59; // @[Parameters.scala 137:67]
  wire [40:0] _T_61; // @[Parameters.scala 137:49]
  wire [40:0] _T_63; // @[Parameters.scala 137:52]
  wire  _T_64; // @[Parameters.scala 137:67]
  wire [39:0] _T_65; // @[Parameters.scala 137:31]
  wire [40:0] _T_66; // @[Parameters.scala 137:49]
  wire [40:0] _T_68; // @[Parameters.scala 137:52]
  wire  _T_69; // @[Parameters.scala 137:67]
  wire [39:0] _T_70; // @[Parameters.scala 137:31]
  wire [40:0] _T_71; // @[Parameters.scala 137:49]
  wire [40:0] _T_73; // @[Parameters.scala 137:52]
  wire  _T_74; // @[Parameters.scala 137:67]
  wire [39:0] _T_75; // @[Parameters.scala 137:31]
  wire [40:0] _T_76; // @[Parameters.scala 137:49]
  wire [40:0] _T_78; // @[Parameters.scala 137:52]
  wire  _T_79; // @[Parameters.scala 137:67]
  wire  _T_81; // @[TLB.scala 195:67]
  wire  _T_82; // @[TLB.scala 195:67]
  wire  _T_83; // @[TLB.scala 195:67]
  wire  _T_84; // @[TLB.scala 195:67]
  wire  _T_85; // @[TLB.scala 195:67]
  wire  legal_address; // @[TLB.scala 195:67]
  wire [40:0] _T_94; // @[Parameters.scala 137:52]
  wire  _T_95; // @[Parameters.scala 137:67]
  wire  cacheable; // @[TLB.scala 197:19]
  wire [39:0] _T_155; // @[Parameters.scala 137:31]
  wire [40:0] _T_156; // @[Parameters.scala 137:49]
  wire [40:0] _T_158; // @[Parameters.scala 137:52]
  wire  _T_159; // @[Parameters.scala 137:67]
  wire [40:0] _T_172; // @[Parameters.scala 137:52]
  wire  _T_173; // @[Parameters.scala 137:67]
  wire  _T_180; // @[TLBPermissions.scala 82:66]
  wire  _T_193; // @[TLB.scala 200:39]
  wire  deny_access_to_debug; // @[TLB.scala 200:48]
  wire  _T_206; // @[TLB.scala 201:41]
  wire  prot_r; // @[TLB.scala 201:66]
  wire [39:0] _T_217; // @[Parameters.scala 137:31]
  wire [40:0] _T_218; // @[Parameters.scala 137:49]
  wire [40:0] _T_220; // @[Parameters.scala 137:52]
  wire  _T_221; // @[Parameters.scala 137:67]
  wire [40:0] _T_225; // @[Parameters.scala 137:52]
  wire  _T_226; // @[Parameters.scala 137:67]
  wire  _T_228; // @[Parameters.scala 549:89]
  wire  _T_229; // @[Parameters.scala 549:89]
  wire  _T_239; // @[TLB.scala 197:19]
  wire  _T_241; // @[TLB.scala 202:45]
  wire  prot_w; // @[TLB.scala 202:70]
  wire  prot_al; // @[TLB.scala 197:19]
  wire [40:0] _T_341; // @[Parameters.scala 137:52]
  wire  _T_342; // @[Parameters.scala 137:67]
  wire  _T_353; // @[Parameters.scala 549:89]
  wire  _T_354; // @[Parameters.scala 549:89]
  wire  _T_370; // @[TLB.scala 197:19]
  wire  _T_372; // @[TLB.scala 206:40]
  wire  prot_x; // @[TLB.scala 206:65]
  wire [40:0] _T_393; // @[Parameters.scala 137:52]
  wire  _T_394; // @[Parameters.scala 137:67]
  wire [40:0] _T_398; // @[Parameters.scala 137:52]
  wire  _T_399; // @[Parameters.scala 137:67]
  wire  _T_410; // @[Parameters.scala 549:89]
  wire  _T_411; // @[Parameters.scala 549:89]
  wire  _T_412; // @[Parameters.scala 549:89]
  wire  prot_eff; // @[TLB.scala 197:19]
  wire  _T_417; // @[package.scala 64:59]
  wire  _T_418; // @[package.scala 64:59]
  wire  _T_419; // @[package.scala 64:59]
  wire [26:0] _T_420; // @[TLB.scala 88:41]
  wire  _T_422; // @[TLB.scala 88:66]
  wire  sector_hits_0; // @[TLB.scala 87:40]
  wire  _T_423; // @[package.scala 64:59]
  wire  _T_424; // @[package.scala 64:59]
  wire  _T_425; // @[package.scala 64:59]
  wire [26:0] _T_426; // @[TLB.scala 88:41]
  wire  _T_428; // @[TLB.scala 88:66]
  wire  sector_hits_1; // @[TLB.scala 87:40]
  wire  _T_429; // @[package.scala 64:59]
  wire  _T_430; // @[package.scala 64:59]
  wire  _T_431; // @[package.scala 64:59]
  wire [26:0] _T_432; // @[TLB.scala 88:41]
  wire  _T_434; // @[TLB.scala 88:66]
  wire  sector_hits_2; // @[TLB.scala 87:40]
  wire  _T_435; // @[package.scala 64:59]
  wire  _T_436; // @[package.scala 64:59]
  wire  _T_437; // @[package.scala 64:59]
  wire [26:0] _T_438; // @[TLB.scala 88:41]
  wire  _T_440; // @[TLB.scala 88:66]
  wire  sector_hits_3; // @[TLB.scala 87:40]
  wire  _T_441; // @[package.scala 64:59]
  wire  _T_442; // @[package.scala 64:59]
  wire  _T_443; // @[package.scala 64:59]
  wire [26:0] _T_444; // @[TLB.scala 88:41]
  wire  _T_446; // @[TLB.scala 88:66]
  wire  sector_hits_4; // @[TLB.scala 87:40]
  wire  _T_447; // @[package.scala 64:59]
  wire  _T_448; // @[package.scala 64:59]
  wire  _T_449; // @[package.scala 64:59]
  wire [26:0] _T_450; // @[TLB.scala 88:41]
  wire  _T_452; // @[TLB.scala 88:66]
  wire  sector_hits_5; // @[TLB.scala 87:40]
  wire  _T_453; // @[package.scala 64:59]
  wire  _T_454; // @[package.scala 64:59]
  wire  _T_455; // @[package.scala 64:59]
  wire [26:0] _T_456; // @[TLB.scala 88:41]
  wire  _T_458; // @[TLB.scala 88:66]
  wire  sector_hits_6; // @[TLB.scala 87:40]
  wire  _T_459; // @[package.scala 64:59]
  wire  _T_460; // @[package.scala 64:59]
  wire  _T_461; // @[package.scala 64:59]
  wire [26:0] _T_462; // @[TLB.scala 88:41]
  wire  _T_464; // @[TLB.scala 88:66]
  wire  sector_hits_7; // @[TLB.scala 87:40]
  wire  _T_469; // @[TLB.scala 95:77]
  wire  _T_471; // @[TLB.scala 95:29]
  wire  _T_472; // @[TLB.scala 94:28]
  wire  _T_476; // @[TLB.scala 95:77]
  wire  _T_477; // @[TLB.scala 95:40]
  wire  superpage_hits_0; // @[TLB.scala 95:29]
  wire  _T_489; // @[TLB.scala 95:77]
  wire  _T_491; // @[TLB.scala 95:29]
  wire  _T_492; // @[TLB.scala 94:28]
  wire  _T_496; // @[TLB.scala 95:77]
  wire  _T_497; // @[TLB.scala 95:40]
  wire  superpage_hits_1; // @[TLB.scala 95:29]
  wire  _T_509; // @[TLB.scala 95:77]
  wire  _T_511; // @[TLB.scala 95:29]
  wire  _T_512; // @[TLB.scala 94:28]
  wire  _T_516; // @[TLB.scala 95:77]
  wire  _T_517; // @[TLB.scala 95:40]
  wire  superpage_hits_2; // @[TLB.scala 95:29]
  wire  _T_529; // @[TLB.scala 95:77]
  wire  _T_531; // @[TLB.scala 95:29]
  wire  _T_532; // @[TLB.scala 94:28]
  wire  _T_536; // @[TLB.scala 95:77]
  wire  _T_537; // @[TLB.scala 95:40]
  wire  superpage_hits_3; // @[TLB.scala 95:29]
  wire  _GEN_1; // @[TLB.scala 100:18]
  wire  _GEN_2; // @[TLB.scala 100:18]
  wire  _GEN_3; // @[TLB.scala 100:18]
  wire  _T_549; // @[TLB.scala 100:18]
  wire  hitsVec_0; // @[TLB.scala 211:44]
  wire  _GEN_5; // @[TLB.scala 100:18]
  wire  _GEN_6; // @[TLB.scala 100:18]
  wire  _GEN_7; // @[TLB.scala 100:18]
  wire  _T_554; // @[TLB.scala 100:18]
  wire  hitsVec_1; // @[TLB.scala 211:44]
  wire  _GEN_9; // @[TLB.scala 100:18]
  wire  _GEN_10; // @[TLB.scala 100:18]
  wire  _GEN_11; // @[TLB.scala 100:18]
  wire  _T_559; // @[TLB.scala 100:18]
  wire  hitsVec_2; // @[TLB.scala 211:44]
  wire  _GEN_13; // @[TLB.scala 100:18]
  wire  _GEN_14; // @[TLB.scala 100:18]
  wire  _GEN_15; // @[TLB.scala 100:18]
  wire  _T_564; // @[TLB.scala 100:18]
  wire  hitsVec_3; // @[TLB.scala 211:44]
  wire  _GEN_17; // @[TLB.scala 100:18]
  wire  _GEN_18; // @[TLB.scala 100:18]
  wire  _GEN_19; // @[TLB.scala 100:18]
  wire  _T_569; // @[TLB.scala 100:18]
  wire  hitsVec_4; // @[TLB.scala 211:44]
  wire  _GEN_21; // @[TLB.scala 100:18]
  wire  _GEN_22; // @[TLB.scala 100:18]
  wire  _GEN_23; // @[TLB.scala 100:18]
  wire  _T_574; // @[TLB.scala 100:18]
  wire  hitsVec_5; // @[TLB.scala 211:44]
  wire  _GEN_25; // @[TLB.scala 100:18]
  wire  _GEN_26; // @[TLB.scala 100:18]
  wire  _GEN_27; // @[TLB.scala 100:18]
  wire  _T_579; // @[TLB.scala 100:18]
  wire  hitsVec_6; // @[TLB.scala 211:44]
  wire  _GEN_29; // @[TLB.scala 100:18]
  wire  _GEN_30; // @[TLB.scala 100:18]
  wire  _GEN_31; // @[TLB.scala 100:18]
  wire  _T_584; // @[TLB.scala 100:18]
  wire  hitsVec_7; // @[TLB.scala 211:44]
  wire  hitsVec_8; // @[TLB.scala 211:44]
  wire  hitsVec_9; // @[TLB.scala 211:44]
  wire  hitsVec_10; // @[TLB.scala 211:44]
  wire  hitsVec_11; // @[TLB.scala 211:44]
  wire  _T_673; // @[TLB.scala 95:77]
  wire  _T_675; // @[TLB.scala 95:29]
  wire  _T_680; // @[TLB.scala 95:77]
  wire  _T_681; // @[TLB.scala 95:40]
  wire  _T_682; // @[TLB.scala 95:29]
  wire  _T_687; // @[TLB.scala 95:77]
  wire  _T_688; // @[TLB.scala 95:40]
  wire  _T_689; // @[TLB.scala 95:29]
  wire  hitsVec_12; // @[TLB.scala 211:44]
  wire [5:0] _T_694; // @[Cat.scala 29:58]
  wire [12:0] real_hits; // @[Cat.scala 29:58]
  wire [13:0] hits; // @[Cat.scala 29:58]
  wire [34:0] _GEN_33;
  wire [34:0] _GEN_34;
  wire [34:0] _GEN_35;
  wire [34:0] _GEN_37;
  wire [34:0] _GEN_38;
  wire [34:0] _GEN_39;
  wire [34:0] _GEN_41;
  wire [34:0] _GEN_42;
  wire [34:0] _GEN_43;
  wire [34:0] _GEN_45;
  wire [34:0] _GEN_46;
  wire [34:0] _GEN_47;
  wire [34:0] _GEN_49;
  wire [34:0] _GEN_50;
  wire [34:0] _GEN_51;
  wire [34:0] _GEN_53;
  wire [34:0] _GEN_54;
  wire [34:0] _GEN_55;
  wire [34:0] _GEN_57;
  wire [34:0] _GEN_58;
  wire [34:0] _GEN_59;
  wire [34:0] _GEN_61;
  wire [34:0] _GEN_62;
  wire [34:0] _GEN_63;
  wire [26:0] _T_876; // @[TLB.scala 109:28]
  wire [26:0] _GEN_985; // @[TLB.scala 109:47]
  wire [26:0] _T_877; // @[TLB.scala 109:47]
  wire [26:0] _T_883; // @[TLB.scala 109:47]
  wire [19:0] _T_885; // @[Cat.scala 29:58]
  wire [26:0] _T_907; // @[TLB.scala 109:28]
  wire [26:0] _GEN_987; // @[TLB.scala 109:47]
  wire [26:0] _T_908; // @[TLB.scala 109:47]
  wire [26:0] _T_914; // @[TLB.scala 109:47]
  wire [19:0] _T_916; // @[Cat.scala 29:58]
  wire [26:0] _T_938; // @[TLB.scala 109:28]
  wire [26:0] _GEN_989; // @[TLB.scala 109:47]
  wire [26:0] _T_939; // @[TLB.scala 109:47]
  wire [26:0] _T_945; // @[TLB.scala 109:47]
  wire [19:0] _T_947; // @[Cat.scala 29:58]
  wire [26:0] _T_969; // @[TLB.scala 109:28]
  wire [26:0] _GEN_991; // @[TLB.scala 109:47]
  wire [26:0] _T_970; // @[TLB.scala 109:47]
  wire [26:0] _T_976; // @[TLB.scala 109:47]
  wire [19:0] _T_978; // @[Cat.scala 29:58]
  wire [26:0] _GEN_993; // @[TLB.scala 109:47]
  wire [26:0] _T_1001; // @[TLB.scala 109:47]
  wire [26:0] _T_1007; // @[TLB.scala 109:47]
  wire [19:0] _T_1009; // @[Cat.scala 29:58]
  wire [19:0] _T_1011; // @[Mux.scala 27:72]
  wire [19:0] _T_1012; // @[Mux.scala 27:72]
  wire [19:0] _T_1013; // @[Mux.scala 27:72]
  wire [19:0] _T_1014; // @[Mux.scala 27:72]
  wire [19:0] _T_1015; // @[Mux.scala 27:72]
  wire [19:0] _T_1016; // @[Mux.scala 27:72]
  wire [19:0] _T_1017; // @[Mux.scala 27:72]
  wire [19:0] _T_1018; // @[Mux.scala 27:72]
  wire [19:0] _T_1019; // @[Mux.scala 27:72]
  wire [19:0] _T_1020; // @[Mux.scala 27:72]
  wire [19:0] _T_1021; // @[Mux.scala 27:72]
  wire [19:0] _T_1022; // @[Mux.scala 27:72]
  wire [19:0] _T_1023; // @[Mux.scala 27:72]
  wire [19:0] _T_1024; // @[Mux.scala 27:72]
  wire [19:0] _T_1025; // @[Mux.scala 27:72]
  wire [19:0] _T_1026; // @[Mux.scala 27:72]
  wire [19:0] _T_1027; // @[Mux.scala 27:72]
  wire [19:0] _T_1028; // @[Mux.scala 27:72]
  wire [19:0] _T_1029; // @[Mux.scala 27:72]
  wire [19:0] _T_1030; // @[Mux.scala 27:72]
  wire [19:0] _T_1031; // @[Mux.scala 27:72]
  wire [19:0] _T_1032; // @[Mux.scala 27:72]
  wire [19:0] _T_1033; // @[Mux.scala 27:72]
  wire [19:0] _T_1034; // @[Mux.scala 27:72]
  wire [19:0] _T_1035; // @[Mux.scala 27:72]
  wire [19:0] _T_1036; // @[Mux.scala 27:72]
  wire [19:0] ppn; // @[Mux.scala 27:72]
  wire  _T_1039; // @[TLB.scala 223:25]
  wire  _T_1041; // @[PTW.scala 69:44]
  wire  _T_1042; // @[PTW.scala 69:38]
  wire  _T_1043; // @[PTW.scala 69:32]
  wire  _T_1044; // @[PTW.scala 69:52]
  wire  _T_1045; // @[PTW.scala 73:35]
  wire  _T_1051; // @[PTW.scala 74:35]
  wire  _T_1052; // @[PTW.scala 74:40]
  wire  _T_1058; // @[PTW.scala 75:35]
  wire [7:0] _T_1068; // @[TLB.scala 123:24]
  wire [34:0] _T_1076; // @[TLB.scala 123:24]
  wire  _GEN_64; // @[TLB.scala 240:34]
  wire  _T_1077; // @[TLB.scala 242:40]
  wire  _T_1078; // @[TLB.scala 243:82]
  wire  _GEN_67; // @[TLB.scala 243:89]
  wire  _T_1095; // @[TLB.scala 243:82]
  wire  _GEN_71; // @[TLB.scala 243:89]
  wire  _T_1112; // @[TLB.scala 243:82]
  wire  _GEN_75; // @[TLB.scala 243:89]
  wire  _T_1129; // @[TLB.scala 243:82]
  wire  _GEN_79; // @[TLB.scala 243:89]
  wire [2:0] _T_1146; // @[TLB.scala 248:22]
  wire  _T_1147; // @[TLB.scala 249:65]
  wire  _GEN_81; // @[TLB.scala 250:32]
  wire  _GEN_82; // @[TLB.scala 250:32]
  wire  _GEN_83; // @[TLB.scala 250:32]
  wire  _GEN_84; // @[TLB.scala 250:32]
  wire  _GEN_995; // @[TLB.scala 122:16]
  wire  _GEN_85; // @[TLB.scala 122:16]
  wire  _GEN_996; // @[TLB.scala 122:16]
  wire  _GEN_86; // @[TLB.scala 122:16]
  wire  _GEN_997; // @[TLB.scala 122:16]
  wire  _GEN_87; // @[TLB.scala 122:16]
  wire  _GEN_998; // @[TLB.scala 122:16]
  wire  _GEN_88; // @[TLB.scala 122:16]
  wire  _GEN_93; // @[TLB.scala 252:34]
  wire  _GEN_94; // @[TLB.scala 252:34]
  wire  _GEN_95; // @[TLB.scala 252:34]
  wire  _GEN_96; // @[TLB.scala 252:34]
  wire  _GEN_97; // @[TLB.scala 249:72]
  wire  _GEN_98; // @[TLB.scala 249:72]
  wire  _GEN_99; // @[TLB.scala 249:72]
  wire  _GEN_100; // @[TLB.scala 249:72]
  wire  _T_1165; // @[TLB.scala 249:65]
  wire  _GEN_107; // @[TLB.scala 250:32]
  wire  _GEN_108; // @[TLB.scala 250:32]
  wire  _GEN_109; // @[TLB.scala 250:32]
  wire  _GEN_110; // @[TLB.scala 250:32]
  wire  _GEN_111; // @[TLB.scala 122:16]
  wire  _GEN_112; // @[TLB.scala 122:16]
  wire  _GEN_113; // @[TLB.scala 122:16]
  wire  _GEN_114; // @[TLB.scala 122:16]
  wire  _GEN_119; // @[TLB.scala 252:34]
  wire  _GEN_120; // @[TLB.scala 252:34]
  wire  _GEN_121; // @[TLB.scala 252:34]
  wire  _GEN_122; // @[TLB.scala 252:34]
  wire  _GEN_123; // @[TLB.scala 249:72]
  wire  _GEN_124; // @[TLB.scala 249:72]
  wire  _GEN_125; // @[TLB.scala 249:72]
  wire  _GEN_126; // @[TLB.scala 249:72]
  wire  _T_1183; // @[TLB.scala 249:65]
  wire  _GEN_133; // @[TLB.scala 250:32]
  wire  _GEN_134; // @[TLB.scala 250:32]
  wire  _GEN_135; // @[TLB.scala 250:32]
  wire  _GEN_136; // @[TLB.scala 250:32]
  wire  _GEN_137; // @[TLB.scala 122:16]
  wire  _GEN_138; // @[TLB.scala 122:16]
  wire  _GEN_139; // @[TLB.scala 122:16]
  wire  _GEN_140; // @[TLB.scala 122:16]
  wire  _GEN_145; // @[TLB.scala 252:34]
  wire  _GEN_146; // @[TLB.scala 252:34]
  wire  _GEN_147; // @[TLB.scala 252:34]
  wire  _GEN_148; // @[TLB.scala 252:34]
  wire  _GEN_149; // @[TLB.scala 249:72]
  wire  _GEN_150; // @[TLB.scala 249:72]
  wire  _GEN_151; // @[TLB.scala 249:72]
  wire  _GEN_152; // @[TLB.scala 249:72]
  wire  _T_1201; // @[TLB.scala 249:65]
  wire  _GEN_159; // @[TLB.scala 250:32]
  wire  _GEN_160; // @[TLB.scala 250:32]
  wire  _GEN_161; // @[TLB.scala 250:32]
  wire  _GEN_162; // @[TLB.scala 250:32]
  wire  _GEN_163; // @[TLB.scala 122:16]
  wire  _GEN_164; // @[TLB.scala 122:16]
  wire  _GEN_165; // @[TLB.scala 122:16]
  wire  _GEN_166; // @[TLB.scala 122:16]
  wire  _GEN_171; // @[TLB.scala 252:34]
  wire  _GEN_172; // @[TLB.scala 252:34]
  wire  _GEN_173; // @[TLB.scala 252:34]
  wire  _GEN_174; // @[TLB.scala 252:34]
  wire  _GEN_175; // @[TLB.scala 249:72]
  wire  _GEN_176; // @[TLB.scala 249:72]
  wire  _GEN_177; // @[TLB.scala 249:72]
  wire  _GEN_178; // @[TLB.scala 249:72]
  wire  _T_1219; // @[TLB.scala 249:65]
  wire  _GEN_185; // @[TLB.scala 250:32]
  wire  _GEN_186; // @[TLB.scala 250:32]
  wire  _GEN_187; // @[TLB.scala 250:32]
  wire  _GEN_188; // @[TLB.scala 250:32]
  wire  _GEN_189; // @[TLB.scala 122:16]
  wire  _GEN_190; // @[TLB.scala 122:16]
  wire  _GEN_191; // @[TLB.scala 122:16]
  wire  _GEN_192; // @[TLB.scala 122:16]
  wire  _GEN_197; // @[TLB.scala 252:34]
  wire  _GEN_198; // @[TLB.scala 252:34]
  wire  _GEN_199; // @[TLB.scala 252:34]
  wire  _GEN_200; // @[TLB.scala 252:34]
  wire  _GEN_201; // @[TLB.scala 249:72]
  wire  _GEN_202; // @[TLB.scala 249:72]
  wire  _GEN_203; // @[TLB.scala 249:72]
  wire  _GEN_204; // @[TLB.scala 249:72]
  wire  _T_1237; // @[TLB.scala 249:65]
  wire  _GEN_211; // @[TLB.scala 250:32]
  wire  _GEN_212; // @[TLB.scala 250:32]
  wire  _GEN_213; // @[TLB.scala 250:32]
  wire  _GEN_214; // @[TLB.scala 250:32]
  wire  _GEN_215; // @[TLB.scala 122:16]
  wire  _GEN_216; // @[TLB.scala 122:16]
  wire  _GEN_217; // @[TLB.scala 122:16]
  wire  _GEN_218; // @[TLB.scala 122:16]
  wire  _GEN_223; // @[TLB.scala 252:34]
  wire  _GEN_224; // @[TLB.scala 252:34]
  wire  _GEN_225; // @[TLB.scala 252:34]
  wire  _GEN_226; // @[TLB.scala 252:34]
  wire  _GEN_227; // @[TLB.scala 249:72]
  wire  _GEN_228; // @[TLB.scala 249:72]
  wire  _GEN_229; // @[TLB.scala 249:72]
  wire  _GEN_230; // @[TLB.scala 249:72]
  wire  _T_1255; // @[TLB.scala 249:65]
  wire  _GEN_237; // @[TLB.scala 250:32]
  wire  _GEN_238; // @[TLB.scala 250:32]
  wire  _GEN_239; // @[TLB.scala 250:32]
  wire  _GEN_240; // @[TLB.scala 250:32]
  wire  _GEN_241; // @[TLB.scala 122:16]
  wire  _GEN_242; // @[TLB.scala 122:16]
  wire  _GEN_243; // @[TLB.scala 122:16]
  wire  _GEN_244; // @[TLB.scala 122:16]
  wire  _GEN_249; // @[TLB.scala 252:34]
  wire  _GEN_250; // @[TLB.scala 252:34]
  wire  _GEN_251; // @[TLB.scala 252:34]
  wire  _GEN_252; // @[TLB.scala 252:34]
  wire  _GEN_253; // @[TLB.scala 249:72]
  wire  _GEN_254; // @[TLB.scala 249:72]
  wire  _GEN_255; // @[TLB.scala 249:72]
  wire  _GEN_256; // @[TLB.scala 249:72]
  wire  _T_1273; // @[TLB.scala 249:65]
  wire  _GEN_263; // @[TLB.scala 250:32]
  wire  _GEN_264; // @[TLB.scala 250:32]
  wire  _GEN_265; // @[TLB.scala 250:32]
  wire  _GEN_266; // @[TLB.scala 250:32]
  wire  _GEN_267; // @[TLB.scala 122:16]
  wire  _GEN_268; // @[TLB.scala 122:16]
  wire  _GEN_269; // @[TLB.scala 122:16]
  wire  _GEN_270; // @[TLB.scala 122:16]
  wire  _GEN_275; // @[TLB.scala 252:34]
  wire  _GEN_276; // @[TLB.scala 252:34]
  wire  _GEN_277; // @[TLB.scala 252:34]
  wire  _GEN_278; // @[TLB.scala 252:34]
  wire  _GEN_279; // @[TLB.scala 249:72]
  wire  _GEN_280; // @[TLB.scala 249:72]
  wire  _GEN_281; // @[TLB.scala 249:72]
  wire  _GEN_282; // @[TLB.scala 249:72]
  wire  _GEN_291; // @[TLB.scala 242:54]
  wire  _GEN_295; // @[TLB.scala 242:54]
  wire  _GEN_299; // @[TLB.scala 242:54]
  wire  _GEN_303; // @[TLB.scala 242:54]
  wire  _GEN_305; // @[TLB.scala 242:54]
  wire  _GEN_306; // @[TLB.scala 242:54]
  wire  _GEN_307; // @[TLB.scala 242:54]
  wire  _GEN_308; // @[TLB.scala 242:54]
  wire  _GEN_315; // @[TLB.scala 242:54]
  wire  _GEN_316; // @[TLB.scala 242:54]
  wire  _GEN_317; // @[TLB.scala 242:54]
  wire  _GEN_318; // @[TLB.scala 242:54]
  wire  _GEN_325; // @[TLB.scala 242:54]
  wire  _GEN_326; // @[TLB.scala 242:54]
  wire  _GEN_327; // @[TLB.scala 242:54]
  wire  _GEN_328; // @[TLB.scala 242:54]
  wire  _GEN_335; // @[TLB.scala 242:54]
  wire  _GEN_336; // @[TLB.scala 242:54]
  wire  _GEN_337; // @[TLB.scala 242:54]
  wire  _GEN_338; // @[TLB.scala 242:54]
  wire  _GEN_345; // @[TLB.scala 242:54]
  wire  _GEN_346; // @[TLB.scala 242:54]
  wire  _GEN_347; // @[TLB.scala 242:54]
  wire  _GEN_348; // @[TLB.scala 242:54]
  wire  _GEN_355; // @[TLB.scala 242:54]
  wire  _GEN_356; // @[TLB.scala 242:54]
  wire  _GEN_357; // @[TLB.scala 242:54]
  wire  _GEN_358; // @[TLB.scala 242:54]
  wire  _GEN_365; // @[TLB.scala 242:54]
  wire  _GEN_366; // @[TLB.scala 242:54]
  wire  _GEN_367; // @[TLB.scala 242:54]
  wire  _GEN_368; // @[TLB.scala 242:54]
  wire  _GEN_375; // @[TLB.scala 242:54]
  wire  _GEN_376; // @[TLB.scala 242:54]
  wire  _GEN_377; // @[TLB.scala 242:54]
  wire  _GEN_378; // @[TLB.scala 242:54]
  wire  _GEN_387; // @[TLB.scala 237:68]
  wire  _GEN_391; // @[TLB.scala 237:68]
  wire  _GEN_395; // @[TLB.scala 237:68]
  wire  _GEN_399; // @[TLB.scala 237:68]
  wire  _GEN_403; // @[TLB.scala 237:68]
  wire  _GEN_405; // @[TLB.scala 237:68]
  wire  _GEN_406; // @[TLB.scala 237:68]
  wire  _GEN_407; // @[TLB.scala 237:68]
  wire  _GEN_408; // @[TLB.scala 237:68]
  wire  _GEN_415; // @[TLB.scala 237:68]
  wire  _GEN_416; // @[TLB.scala 237:68]
  wire  _GEN_417; // @[TLB.scala 237:68]
  wire  _GEN_418; // @[TLB.scala 237:68]
  wire  _GEN_425; // @[TLB.scala 237:68]
  wire  _GEN_426; // @[TLB.scala 237:68]
  wire  _GEN_427; // @[TLB.scala 237:68]
  wire  _GEN_428; // @[TLB.scala 237:68]
  wire  _GEN_435; // @[TLB.scala 237:68]
  wire  _GEN_436; // @[TLB.scala 237:68]
  wire  _GEN_437; // @[TLB.scala 237:68]
  wire  _GEN_438; // @[TLB.scala 237:68]
  wire  _GEN_445; // @[TLB.scala 237:68]
  wire  _GEN_446; // @[TLB.scala 237:68]
  wire  _GEN_447; // @[TLB.scala 237:68]
  wire  _GEN_448; // @[TLB.scala 237:68]
  wire  _GEN_455; // @[TLB.scala 237:68]
  wire  _GEN_456; // @[TLB.scala 237:68]
  wire  _GEN_457; // @[TLB.scala 237:68]
  wire  _GEN_458; // @[TLB.scala 237:68]
  wire  _GEN_465; // @[TLB.scala 237:68]
  wire  _GEN_466; // @[TLB.scala 237:68]
  wire  _GEN_467; // @[TLB.scala 237:68]
  wire  _GEN_468; // @[TLB.scala 237:68]
  wire  _GEN_475; // @[TLB.scala 237:68]
  wire  _GEN_476; // @[TLB.scala 237:68]
  wire  _GEN_477; // @[TLB.scala 237:68]
  wire  _GEN_478; // @[TLB.scala 237:68]
  wire  _GEN_487; // @[TLB.scala 217:20]
  wire  _GEN_491; // @[TLB.scala 217:20]
  wire  _GEN_495; // @[TLB.scala 217:20]
  wire  _GEN_499; // @[TLB.scala 217:20]
  wire  _GEN_503; // @[TLB.scala 217:20]
  wire  _GEN_505; // @[TLB.scala 217:20]
  wire  _GEN_506; // @[TLB.scala 217:20]
  wire  _GEN_507; // @[TLB.scala 217:20]
  wire  _GEN_508; // @[TLB.scala 217:20]
  wire  _GEN_515; // @[TLB.scala 217:20]
  wire  _GEN_516; // @[TLB.scala 217:20]
  wire  _GEN_517; // @[TLB.scala 217:20]
  wire  _GEN_518; // @[TLB.scala 217:20]
  wire  _GEN_525; // @[TLB.scala 217:20]
  wire  _GEN_526; // @[TLB.scala 217:20]
  wire  _GEN_527; // @[TLB.scala 217:20]
  wire  _GEN_528; // @[TLB.scala 217:20]
  wire  _GEN_535; // @[TLB.scala 217:20]
  wire  _GEN_536; // @[TLB.scala 217:20]
  wire  _GEN_537; // @[TLB.scala 217:20]
  wire  _GEN_538; // @[TLB.scala 217:20]
  wire  _GEN_545; // @[TLB.scala 217:20]
  wire  _GEN_546; // @[TLB.scala 217:20]
  wire  _GEN_547; // @[TLB.scala 217:20]
  wire  _GEN_548; // @[TLB.scala 217:20]
  wire  _GEN_555; // @[TLB.scala 217:20]
  wire  _GEN_556; // @[TLB.scala 217:20]
  wire  _GEN_557; // @[TLB.scala 217:20]
  wire  _GEN_558; // @[TLB.scala 217:20]
  wire  _GEN_565; // @[TLB.scala 217:20]
  wire  _GEN_566; // @[TLB.scala 217:20]
  wire  _GEN_567; // @[TLB.scala 217:20]
  wire  _GEN_568; // @[TLB.scala 217:20]
  wire  _GEN_575; // @[TLB.scala 217:20]
  wire  _GEN_576; // @[TLB.scala 217:20]
  wire  _GEN_577; // @[TLB.scala 217:20]
  wire  _GEN_578; // @[TLB.scala 217:20]
  wire [5:0] _T_1761; // @[Cat.scala 29:58]
  wire [13:0] ptw_ae_array; // @[Cat.scala 29:58]
  wire [5:0] _T_1775; // @[Cat.scala 29:58]
  wire [12:0] _T_1782; // @[Cat.scala 29:58]
  wire [12:0] priv_x_ok; // @[TLB.scala 262:22]
  wire [5:0] _T_1839; // @[Cat.scala 29:58]
  wire [12:0] _T_1846; // @[Cat.scala 29:58]
  wire [12:0] _T_1875; // @[TLB.scala 265:39]
  wire [13:0] x_array; // @[Cat.scala 29:58]
  wire [1:0] _T_1907; // @[Bitwise.scala 72:12]
  wire [5:0] _T_1912; // @[Cat.scala 29:58]
  wire [13:0] _T_1919; // @[Cat.scala 29:58]
  wire [13:0] px_array; // @[TLB.scala 268:87]
  wire [1:0] _T_1935; // @[Bitwise.scala 72:12]
  wire [5:0] _T_1940; // @[Cat.scala 29:58]
  wire [13:0] c_array; // @[Cat.scala 29:58]
  wire [39:0] _T_2005; // @[TLB.scala 285:43]
  wire  _T_2007; // @[TLB.scala 286:61]
  wire  _T_2008; // @[TLB.scala 286:82]
  wire  _T_2009; // @[TLB.scala 286:67]
  wire  bad_va; // @[TLB.scala 280:117]
  wire [13:0] _T_2112; // @[TLB.scala 318:33]
  wire [13:0] pf_inst_array; // @[TLB.scala 318:23]
  wire  tlb_hit; // @[TLB.scala 320:27]
  wire  _T_2114; // @[TLB.scala 321:29]
  wire  tlb_miss; // @[TLB.scala 321:40]
  reg [6:0] _T_2116; // @[Replacement.scala 158:30]
  reg [31:0] _RAND_98;
  reg [2:0] _T_2117; // @[Replacement.scala 158:30]
  reg [31:0] _RAND_99;
  wire  _T_2118; // @[TLB.scala 325:22]
  wire  _T_2119; // @[package.scala 64:59]
  wire  _T_2120; // @[package.scala 64:59]
  wire  _T_2121; // @[package.scala 64:59]
  wire  _T_2122; // @[package.scala 64:59]
  wire  _T_2123; // @[package.scala 64:59]
  wire  _T_2124; // @[package.scala 64:59]
  wire  _T_2125; // @[package.scala 64:59]
  wire [7:0] _T_2132; // @[Cat.scala 29:58]
  wire  _T_2135; // @[OneHot.scala 32:14]
  wire [3:0] _T_2136; // @[OneHot.scala 32:28]
  wire  _T_2139; // @[OneHot.scala 32:14]
  wire [1:0] _T_2140; // @[OneHot.scala 32:28]
  wire [2:0] _T_2143; // @[Cat.scala 29:58]
  wire  _T_2157; // @[Replacement.scala 193:16]
  wire  _T_2161; // @[Replacement.scala 196:16]
  wire [2:0] _T_2163; // @[Cat.scala 29:58]
  wire [2:0] _T_2164; // @[Replacement.scala 193:16]
  wire  _T_2173; // @[Replacement.scala 193:16]
  wire  _T_2177; // @[Replacement.scala 196:16]
  wire [2:0] _T_2179; // @[Cat.scala 29:58]
  wire [2:0] _T_2180; // @[Replacement.scala 196:16]
  wire [6:0] _T_2182; // @[Cat.scala 29:58]
  wire  _T_2183; // @[package.scala 64:59]
  wire  _T_2184; // @[package.scala 64:59]
  wire  _T_2185; // @[package.scala 64:59]
  wire [3:0] _T_2188; // @[Cat.scala 29:58]
  wire  _T_2191; // @[OneHot.scala 32:14]
  wire [1:0] _T_2192; // @[OneHot.scala 32:28]
  wire [1:0] _T_2194; // @[Cat.scala 29:58]
  wire  _T_2203; // @[Replacement.scala 193:16]
  wire  _T_2207; // @[Replacement.scala 196:16]
  wire [2:0] _T_2209; // @[Cat.scala 29:58]
  wire  _T_2219; // @[Misc.scala 182:16]
  wire  _T_2221; // @[Misc.scala 182:61]
  wire  _T_2223; // @[Misc.scala 182:16]
  wire  _T_2225; // @[Misc.scala 182:61]
  wire  _T_2226; // @[Misc.scala 182:49]
  wire  _T_2235; // @[Misc.scala 182:16]
  wire  _T_2237; // @[Misc.scala 182:61]
  wire  _T_2239; // @[Misc.scala 182:16]
  wire  _T_2241; // @[Misc.scala 182:61]
  wire  _T_2242; // @[Misc.scala 182:49]
  wire  _T_2243; // @[Misc.scala 182:16]
  wire  _T_2244; // @[Misc.scala 182:37]
  wire  _T_2245; // @[Misc.scala 182:61]
  wire  _T_2246; // @[Misc.scala 182:49]
  wire  _T_2256; // @[Misc.scala 182:16]
  wire  _T_2258; // @[Misc.scala 182:61]
  wire  _T_2260; // @[Misc.scala 182:16]
  wire  _T_2262; // @[Misc.scala 182:61]
  wire  _T_2263; // @[Misc.scala 182:49]
  wire  _T_2270; // @[Misc.scala 182:16]
  wire  _T_2272; // @[Misc.scala 182:61]
  wire  _T_2279; // @[Misc.scala 182:16]
  wire  _T_2281; // @[Misc.scala 182:61]
  wire  _T_2283; // @[Misc.scala 182:16]
  wire  _T_2284; // @[Misc.scala 182:37]
  wire  _T_2285; // @[Misc.scala 182:61]
  wire  _T_2286; // @[Misc.scala 182:49]
  wire  _T_2287; // @[Misc.scala 182:16]
  wire  _T_2288; // @[Misc.scala 182:37]
  wire  _T_2289; // @[Misc.scala 182:61]
  wire  _T_2290; // @[Misc.scala 182:49]
  wire  _T_2292; // @[Misc.scala 182:37]
  wire  _T_2293; // @[Misc.scala 182:61]
  wire  multipleHits; // @[Misc.scala 182:49]
  wire [13:0] _T_2303; // @[TLB.scala 340:47]
  wire  _T_2304; // @[TLB.scala 340:55]
  wire [13:0] _T_2311; // @[TLB.scala 343:33]
  wire [13:0] _T_2317; // @[TLB.scala 347:33]
  wire  _T_2324; // @[TLB.scala 350:29]
  wire  _T_2330; // @[Decoupled.scala 40:37]
  wire  _T_2331; // @[TLB.scala 359:25]
  wire  _T_2337; // @[Replacement.scala 240:16]
  wire [1:0] _T_2338; // @[Cat.scala 29:58]
  wire [3:0] _T_2341; // @[Cat.scala 29:58]
  wire  _T_2342; // @[TLB.scala 407:16]
  wire  _T_2344; // @[OneHot.scala 47:40]
  wire  _T_2345; // @[OneHot.scala 47:40]
  wire  _T_2346; // @[OneHot.scala 47:40]
  wire  _T_2360; // @[Replacement.scala 240:16]
  wire [1:0] _T_2361; // @[Cat.scala 29:58]
  wire  _T_2367; // @[Replacement.scala 240:16]
  wire [1:0] _T_2368; // @[Cat.scala 29:58]
  wire [1:0] _T_2369; // @[Replacement.scala 240:16]
  wire [2:0] _T_2370; // @[Cat.scala 29:58]
  wire [7:0] _T_2401; // @[Cat.scala 29:58]
  wire  _T_2402; // @[TLB.scala 407:16]
  wire  _T_2404; // @[OneHot.scala 47:40]
  wire  _T_2405; // @[OneHot.scala 47:40]
  wire  _T_2406; // @[OneHot.scala 47:40]
  wire  _T_2407; // @[OneHot.scala 47:40]
  wire  _T_2408; // @[OneHot.scala 47:40]
  wire  _T_2409; // @[OneHot.scala 47:40]
  wire  _T_2410; // @[OneHot.scala 47:40]
  wire  _T_2447; // @[TLB.scala 373:17]
  wire  _T_2448; // @[TLB.scala 373:28]
  wire  _T_2451; // @[TLB.scala 381:72]
  wire  _T_2452; // @[TLB.scala 381:34]
  wire  _T_2454; // @[TLB.scala 381:13]
  wire  _T_2462; // @[TLB.scala 135:61]
  wire  _GEN_681; // @[TLB.scala 143:19]
  wire  _GEN_682; // @[TLB.scala 143:19]
  wire  _GEN_683; // @[TLB.scala 143:19]
  wire  _GEN_684; // @[TLB.scala 143:19]
  wire  _GEN_685; // @[TLB.scala 384:40]
  wire  _GEN_686; // @[TLB.scala 384:40]
  wire  _GEN_687; // @[TLB.scala 384:40]
  wire  _GEN_688; // @[TLB.scala 384:40]
  wire  _T_2617; // @[TLB.scala 135:61]
  wire  _GEN_709; // @[TLB.scala 143:19]
  wire  _GEN_710; // @[TLB.scala 143:19]
  wire  _GEN_711; // @[TLB.scala 143:19]
  wire  _GEN_712; // @[TLB.scala 143:19]
  wire  _GEN_713; // @[TLB.scala 384:40]
  wire  _GEN_714; // @[TLB.scala 384:40]
  wire  _GEN_715; // @[TLB.scala 384:40]
  wire  _GEN_716; // @[TLB.scala 384:40]
  wire  _T_2772; // @[TLB.scala 135:61]
  wire  _GEN_737; // @[TLB.scala 143:19]
  wire  _GEN_738; // @[TLB.scala 143:19]
  wire  _GEN_739; // @[TLB.scala 143:19]
  wire  _GEN_740; // @[TLB.scala 143:19]
  wire  _GEN_741; // @[TLB.scala 384:40]
  wire  _GEN_742; // @[TLB.scala 384:40]
  wire  _GEN_743; // @[TLB.scala 384:40]
  wire  _GEN_744; // @[TLB.scala 384:40]
  wire  _T_2927; // @[TLB.scala 135:61]
  wire  _GEN_765; // @[TLB.scala 143:19]
  wire  _GEN_766; // @[TLB.scala 143:19]
  wire  _GEN_767; // @[TLB.scala 143:19]
  wire  _GEN_768; // @[TLB.scala 143:19]
  wire  _GEN_769; // @[TLB.scala 384:40]
  wire  _GEN_770; // @[TLB.scala 384:40]
  wire  _GEN_771; // @[TLB.scala 384:40]
  wire  _GEN_772; // @[TLB.scala 384:40]
  wire  _T_3082; // @[TLB.scala 135:61]
  wire  _GEN_793; // @[TLB.scala 143:19]
  wire  _GEN_794; // @[TLB.scala 143:19]
  wire  _GEN_795; // @[TLB.scala 143:19]
  wire  _GEN_796; // @[TLB.scala 143:19]
  wire  _GEN_797; // @[TLB.scala 384:40]
  wire  _GEN_798; // @[TLB.scala 384:40]
  wire  _GEN_799; // @[TLB.scala 384:40]
  wire  _GEN_800; // @[TLB.scala 384:40]
  wire  _T_3237; // @[TLB.scala 135:61]
  wire  _GEN_821; // @[TLB.scala 143:19]
  wire  _GEN_822; // @[TLB.scala 143:19]
  wire  _GEN_823; // @[TLB.scala 143:19]
  wire  _GEN_824; // @[TLB.scala 143:19]
  wire  _GEN_825; // @[TLB.scala 384:40]
  wire  _GEN_826; // @[TLB.scala 384:40]
  wire  _GEN_827; // @[TLB.scala 384:40]
  wire  _GEN_828; // @[TLB.scala 384:40]
  wire  _T_3392; // @[TLB.scala 135:61]
  wire  _GEN_849; // @[TLB.scala 143:19]
  wire  _GEN_850; // @[TLB.scala 143:19]
  wire  _GEN_851; // @[TLB.scala 143:19]
  wire  _GEN_852; // @[TLB.scala 143:19]
  wire  _GEN_853; // @[TLB.scala 384:40]
  wire  _GEN_854; // @[TLB.scala 384:40]
  wire  _GEN_855; // @[TLB.scala 384:40]
  wire  _GEN_856; // @[TLB.scala 384:40]
  wire  _T_3547; // @[TLB.scala 135:61]
  wire  _GEN_877; // @[TLB.scala 143:19]
  wire  _GEN_878; // @[TLB.scala 143:19]
  wire  _GEN_879; // @[TLB.scala 143:19]
  wire  _GEN_880; // @[TLB.scala 143:19]
  wire  _GEN_881; // @[TLB.scala 384:40]
  wire  _GEN_882; // @[TLB.scala 384:40]
  wire  _GEN_883; // @[TLB.scala 384:40]
  wire  _GEN_884; // @[TLB.scala 384:40]
  wire  _GEN_890; // @[TLB.scala 143:19]
  wire  _GEN_891; // @[TLB.scala 384:40]
  wire  _GEN_894; // @[TLB.scala 143:19]
  wire  _GEN_895; // @[TLB.scala 384:40]
  wire  _GEN_898; // @[TLB.scala 143:19]
  wire  _GEN_899; // @[TLB.scala 384:40]
  wire  _GEN_902; // @[TLB.scala 143:19]
  wire  _GEN_903; // @[TLB.scala 384:40]
  wire  _GEN_906; // @[TLB.scala 143:19]
  wire  _GEN_907; // @[TLB.scala 384:40]
  wire  _T_3897; // @[TLB.scala 388:24]
  reg [19:0] TLB_1_state; // @[Register tracking TLB_1 state]
  reg [31:0] _RAND_100;
  reg  TLB_1_cov [0:1048575]; // @[Coverage map for TLB_1]
  reg [31:0] _RAND_101;
  wire  TLB_1_cov_read_data; // @[Coverage map for TLB_1]
  wire [19:0] TLB_1_cov_read_addr; // @[Coverage map for TLB_1]
  wire  TLB_1_cov_write_data; // @[Coverage map for TLB_1]
  wire [19:0] TLB_1_cov_write_addr; // @[Coverage map for TLB_1]
  wire  TLB_1_cov_write_mask; // @[Coverage map for TLB_1]
  wire  TLB_1_cov_write_en; // @[Coverage map for TLB_1]
  reg [29:0] TLB_1_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_102;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire  mux_cond_6;
  wire  mux_cond_7;
  wire  mux_cond_8;
  wire  mux_cond_9;
  wire  mux_cond_10;
  wire  mux_cond_11;
  wire  mux_cond_12;
  wire  mux_cond_13;
  wire  mux_cond_14;
  wire  mux_cond_15;
  wire  mux_cond_16;
  wire  mux_cond_17;
  wire  mux_cond_18;
  wire  mux_cond_19;
  wire  mux_cond_20;
  wire  mux_cond_21;
  wire  mux_cond_22;
  wire  mux_cond_23;
  wire  mux_cond_24;
  wire  mux_cond_25;
  wire  mux_cond_26;
  wire  mux_cond_27;
  wire  mux_cond_28;
  wire  mux_cond_29;
  wire  mux_cond_30;
  wire  mux_cond_31;
  wire  mux_cond_32;
  wire  mux_cond_33;
  wire  mux_cond_34;
  wire  mux_cond_35;
  wire  mux_cond_36;
  wire  mux_cond_37;
  wire  mux_cond_38;
  wire  mux_cond_39;
  wire  mux_cond_40;
  wire  mux_cond_41;
  wire  mux_cond_42;
  wire  mux_cond_43;
  wire  mux_cond_44;
  wire  mux_cond_45;
  wire  mux_cond_46;
  wire  mux_cond_47;
  wire  mux_cond_48;
  wire  mux_cond_49;
  wire  mux_cond_50;
  wire  mux_cond_51;
  wire  mux_cond_52;
  wire  mux_cond_53;
  wire  mux_cond_54;
  wire  mux_cond_55;
  wire  mux_cond_56;
  wire  mux_cond_57;
  wire  mux_cond_58;
  wire  mux_cond_59;
  wire  mux_cond_60;
  wire  mux_cond_61;
  wire  mux_cond_62;
  wire  mux_cond_63;
  wire  mux_cond_64;
  wire  mux_cond_65;
  wire  mux_cond_66;
  wire  mux_cond_67;
  wire  mux_cond_68;
  wire [3:0] state_shl;
  wire [19:0] state_pad;
  wire [2:0] r_sectored_repl_addr_shl;
  wire [19:0] r_sectored_repl_addr_pad;
  wire [15:0] r_superpage_repl_addr_shl;
  wire [19:0] r_superpage_repl_addr_pad;
  wire [3:0] r_sectored_hit_addr_shl;
  wire [19:0] r_sectored_hit_addr_pad;
  wire [18:0] special_entry_valid_0_shl;
  wire [19:0] special_entry_valid_0_pad;
  wire [4:0] r_sectored_hit_shl;
  wire [19:0] r_sectored_hit_pad;
  wire [12:0] special_entry_level_shl;
  wire [19:0] special_entry_level_pad;
  wire [18:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [8:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [3:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [18:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [9:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [12:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [12:0] mux_cond_6_shl;
  wire [19:0] mux_cond_6_pad;
  wire [6:0] mux_cond_7_shl;
  wire [19:0] mux_cond_7_pad;
  wire [1:0] mux_cond_8_shl;
  wire [19:0] mux_cond_8_pad;
  wire [17:0] mux_cond_9_shl;
  wire [19:0] mux_cond_9_pad;
  wire [5:0] mux_cond_10_shl;
  wire [19:0] mux_cond_10_pad;
  wire  mux_cond_11_shl;
  wire [19:0] mux_cond_11_pad;
  wire [12:0] mux_cond_12_shl;
  wire [19:0] mux_cond_12_pad;
  wire [15:0] mux_cond_13_shl;
  wire [19:0] mux_cond_13_pad;
  wire [17:0] mux_cond_14_shl;
  wire [19:0] mux_cond_14_pad;
  wire [13:0] mux_cond_15_shl;
  wire [19:0] mux_cond_15_pad;
  wire [18:0] mux_cond_16_shl;
  wire [19:0] mux_cond_16_pad;
  wire [4:0] mux_cond_17_shl;
  wire [19:0] mux_cond_17_pad;
  wire [4:0] mux_cond_18_shl;
  wire [19:0] mux_cond_18_pad;
  wire [19:0] mux_cond_19_shl;
  wire [19:0] mux_cond_19_pad;
  wire [12:0] mux_cond_20_shl;
  wire [19:0] mux_cond_20_pad;
  wire [6:0] mux_cond_21_shl;
  wire [19:0] mux_cond_21_pad;
  wire [11:0] mux_cond_22_shl;
  wire [19:0] mux_cond_22_pad;
  wire  mux_cond_23_shl;
  wire [19:0] mux_cond_23_pad;
  wire  mux_cond_24_shl;
  wire [19:0] mux_cond_24_pad;
  wire [16:0] mux_cond_25_shl;
  wire [19:0] mux_cond_25_pad;
  wire [16:0] mux_cond_26_shl;
  wire [19:0] mux_cond_26_pad;
  wire [4:0] mux_cond_27_shl;
  wire [19:0] mux_cond_27_pad;
  wire [16:0] mux_cond_28_shl;
  wire [19:0] mux_cond_28_pad;
  wire [5:0] mux_cond_29_shl;
  wire [19:0] mux_cond_29_pad;
  wire [11:0] mux_cond_30_shl;
  wire [19:0] mux_cond_30_pad;
  wire [18:0] mux_cond_31_shl;
  wire [19:0] mux_cond_31_pad;
  wire [2:0] mux_cond_32_shl;
  wire [19:0] mux_cond_32_pad;
  wire [15:0] mux_cond_33_shl;
  wire [19:0] mux_cond_33_pad;
  wire [15:0] mux_cond_34_shl;
  wire [19:0] mux_cond_34_pad;
  wire [7:0] mux_cond_35_shl;
  wire [19:0] mux_cond_35_pad;
  wire [9:0] mux_cond_36_shl;
  wire [19:0] mux_cond_36_pad;
  wire [15:0] mux_cond_37_shl;
  wire [19:0] mux_cond_37_pad;
  wire  mux_cond_38_shl;
  wire [19:0] mux_cond_38_pad;
  wire [12:0] mux_cond_39_shl;
  wire [19:0] mux_cond_39_pad;
  wire [15:0] mux_cond_40_shl;
  wire [19:0] mux_cond_40_pad;
  wire [13:0] mux_cond_41_shl;
  wire [19:0] mux_cond_41_pad;
  wire [7:0] mux_cond_42_shl;
  wire [19:0] mux_cond_42_pad;
  wire [2:0] mux_cond_43_shl;
  wire [19:0] mux_cond_43_pad;
  wire [6:0] mux_cond_44_shl;
  wire [19:0] mux_cond_44_pad;
  wire [8:0] mux_cond_45_shl;
  wire [19:0] mux_cond_45_pad;
  wire [13:0] mux_cond_46_shl;
  wire [19:0] mux_cond_46_pad;
  wire [19:0] mux_cond_47_shl;
  wire [19:0] mux_cond_47_pad;
  wire [10:0] mux_cond_48_shl;
  wire [19:0] mux_cond_48_pad;
  wire [2:0] mux_cond_49_shl;
  wire [19:0] mux_cond_49_pad;
  wire [6:0] mux_cond_50_shl;
  wire [19:0] mux_cond_50_pad;
  wire [2:0] mux_cond_51_shl;
  wire [19:0] mux_cond_51_pad;
  wire [8:0] mux_cond_52_shl;
  wire [19:0] mux_cond_52_pad;
  wire [11:0] mux_cond_53_shl;
  wire [19:0] mux_cond_53_pad;
  wire [8:0] mux_cond_54_shl;
  wire [19:0] mux_cond_54_pad;
  wire [12:0] mux_cond_55_shl;
  wire [19:0] mux_cond_55_pad;
  wire [10:0] mux_cond_56_shl;
  wire [19:0] mux_cond_56_pad;
  wire [3:0] mux_cond_57_shl;
  wire [19:0] mux_cond_57_pad;
  wire  mux_cond_58_shl;
  wire [19:0] mux_cond_58_pad;
  wire [11:0] mux_cond_59_shl;
  wire [19:0] mux_cond_59_pad;
  wire [3:0] mux_cond_60_shl;
  wire [19:0] mux_cond_60_pad;
  wire [13:0] mux_cond_61_shl;
  wire [19:0] mux_cond_61_pad;
  wire [8:0] mux_cond_62_shl;
  wire [19:0] mux_cond_62_pad;
  wire  mux_cond_63_shl;
  wire [19:0] mux_cond_63_pad;
  wire [6:0] mux_cond_64_shl;
  wire [19:0] mux_cond_64_pad;
  wire [13:0] mux_cond_65_shl;
  wire [19:0] mux_cond_65_pad;
  wire [4:0] mux_cond_66_shl;
  wire [19:0] mux_cond_66_pad;
  wire [10:0] mux_cond_67_shl;
  wire [19:0] mux_cond_67_pad;
  wire [15:0] mux_cond_68_shl;
  wire [19:0] mux_cond_68_pad;
  wire [17:0] superpage_entries_2_level_shl;
  wire [19:0] superpage_entries_2_level_pad;
  wire [14:0] sectored_entries_7_valid_3_shl;
  wire [19:0] sectored_entries_7_valid_3_pad;
  wire [17:0] superpage_entries_1_level_shl;
  wire [19:0] superpage_entries_1_level_pad;
  wire [11:0] superpage_entries_1_valid_0_shl;
  wire [19:0] superpage_entries_1_valid_0_pad;
  wire [18:0] sectored_entries_3_valid_0_shl;
  wire [19:0] sectored_entries_3_valid_0_pad;
  wire [14:0] sectored_entries_1_valid_3_shl;
  wire [19:0] sectored_entries_1_valid_3_pad;
  wire [14:0] sectored_entries_6_valid_3_shl;
  wire [19:0] sectored_entries_6_valid_3_pad;
  wire [18:0] sectored_entries_1_valid_0_shl;
  wire [19:0] sectored_entries_1_valid_0_pad;
  wire [18:0] sectored_entries_2_valid_0_shl;
  wire [19:0] sectored_entries_2_valid_0_pad;
  wire [14:0] sectored_entries_3_valid_1_shl;
  wire [19:0] sectored_entries_3_valid_1_pad;
  wire [14:0] sectored_entries_5_valid_3_shl;
  wire [19:0] sectored_entries_5_valid_3_pad;
  wire [11:0] superpage_entries_3_valid_0_shl;
  wire [19:0] superpage_entries_3_valid_0_pad;
  wire [14:0] sectored_entries_5_valid_1_shl;
  wire [19:0] sectored_entries_5_valid_1_pad;
  wire [14:0] sectored_entries_0_valid_3_shl;
  wire [19:0] sectored_entries_0_valid_3_pad;
  wire [18:0] sectored_entries_6_valid_0_shl;
  wire [19:0] sectored_entries_6_valid_0_pad;
  wire [18:0] sectored_entries_0_valid_0_shl;
  wire [19:0] sectored_entries_0_valid_0_pad;
  wire [16:0] sectored_entries_4_valid_2_shl;
  wire [19:0] sectored_entries_4_valid_2_pad;
  wire [11:0] superpage_entries_2_valid_0_shl;
  wire [19:0] superpage_entries_2_valid_0_pad;
  wire [14:0] sectored_entries_2_valid_1_shl;
  wire [19:0] sectored_entries_2_valid_1_pad;
  wire [17:0] superpage_entries_0_level_shl;
  wire [19:0] superpage_entries_0_level_pad;
  wire [14:0] sectored_entries_1_valid_1_shl;
  wire [19:0] sectored_entries_1_valid_1_pad;
  wire [14:0] sectored_entries_4_valid_3_shl;
  wire [19:0] sectored_entries_4_valid_3_pad;
  wire [14:0] sectored_entries_0_valid_1_shl;
  wire [19:0] sectored_entries_0_valid_1_pad;
  wire [18:0] sectored_entries_4_valid_0_shl;
  wire [19:0] sectored_entries_4_valid_0_pad;
  wire [16:0] sectored_entries_0_valid_2_shl;
  wire [19:0] sectored_entries_0_valid_2_pad;
  wire [16:0] sectored_entries_1_valid_2_shl;
  wire [19:0] sectored_entries_1_valid_2_pad;
  wire [16:0] sectored_entries_2_valid_2_shl;
  wire [19:0] sectored_entries_2_valid_2_pad;
  wire [18:0] sectored_entries_7_valid_0_shl;
  wire [19:0] sectored_entries_7_valid_0_pad;
  wire [16:0] sectored_entries_5_valid_2_shl;
  wire [19:0] sectored_entries_5_valid_2_pad;
  wire [16:0] sectored_entries_7_valid_2_shl;
  wire [19:0] sectored_entries_7_valid_2_pad;
  wire [14:0] sectored_entries_4_valid_1_shl;
  wire [19:0] sectored_entries_4_valid_1_pad;
  wire [18:0] sectored_entries_5_valid_0_shl;
  wire [19:0] sectored_entries_5_valid_0_pad;
  wire [14:0] sectored_entries_7_valid_1_shl;
  wire [19:0] sectored_entries_7_valid_1_pad;
  wire [17:0] superpage_entries_3_level_shl;
  wire [19:0] superpage_entries_3_level_pad;
  wire [14:0] sectored_entries_3_valid_3_shl;
  wire [19:0] sectored_entries_3_valid_3_pad;
  wire [14:0] sectored_entries_2_valid_3_shl;
  wire [19:0] sectored_entries_2_valid_3_pad;
  wire [11:0] superpage_entries_0_valid_0_shl;
  wire [19:0] superpage_entries_0_valid_0_pad;
  wire [14:0] sectored_entries_6_valid_1_shl;
  wire [19:0] sectored_entries_6_valid_1_pad;
  wire [16:0] sectored_entries_3_valid_2_shl;
  wire [19:0] sectored_entries_3_valid_2_pad;
  wire [16:0] sectored_entries_6_valid_2_shl;
  wire [19:0] sectored_entries_6_valid_2_pad;
  wire [19:0] TLB_1_xor64;
  wire [19:0] TLB_1_xor31;
  wire [19:0] TLB_1_xor65;
  wire [19:0] TLB_1_xor66;
  wire [19:0] TLB_1_xor32;
  wire [19:0] TLB_1_xor15;
  wire [19:0] TLB_1_xor68;
  wire [19:0] TLB_1_xor33;
  wire [19:0] TLB_1_xor69;
  wire [19:0] TLB_1_xor70;
  wire [19:0] TLB_1_xor34;
  wire [19:0] TLB_1_xor16;
  wire [19:0] TLB_1_xor7;
  wire [19:0] TLB_1_xor72;
  wire [19:0] TLB_1_xor35;
  wire [19:0] TLB_1_xor73;
  wire [19:0] TLB_1_xor74;
  wire [19:0] TLB_1_xor36;
  wire [19:0] TLB_1_xor17;
  wire [19:0] TLB_1_xor75;
  wire [19:0] TLB_1_xor76;
  wire [19:0] TLB_1_xor37;
  wire [19:0] TLB_1_xor77;
  wire [19:0] TLB_1_xor78;
  wire [19:0] TLB_1_xor38;
  wire [19:0] TLB_1_xor18;
  wire [19:0] TLB_1_xor8;
  wire [19:0] TLB_1_xor3;
  wire [19:0] TLB_1_xor80;
  wire [19:0] TLB_1_xor39;
  wire [19:0] TLB_1_xor81;
  wire [19:0] TLB_1_xor82;
  wire [19:0] TLB_1_xor40;
  wire [19:0] TLB_1_xor19;
  wire [19:0] TLB_1_xor84;
  wire [19:0] TLB_1_xor41;
  wire [19:0] TLB_1_xor85;
  wire [19:0] TLB_1_xor86;
  wire [19:0] TLB_1_xor42;
  wire [19:0] TLB_1_xor20;
  wire [19:0] TLB_1_xor9;
  wire [19:0] TLB_1_xor88;
  wire [19:0] TLB_1_xor43;
  wire [19:0] TLB_1_xor89;
  wire [19:0] TLB_1_xor90;
  wire [19:0] TLB_1_xor44;
  wire [19:0] TLB_1_xor21;
  wire [19:0] TLB_1_xor91;
  wire [19:0] TLB_1_xor92;
  wire [19:0] TLB_1_xor45;
  wire [19:0] TLB_1_xor93;
  wire [19:0] TLB_1_xor94;
  wire [19:0] TLB_1_xor46;
  wire [19:0] TLB_1_xor22;
  wire [19:0] TLB_1_xor10;
  wire [19:0] TLB_1_xor4;
  wire [19:0] TLB_1_xor1;
  wire [19:0] TLB_1_xor96;
  wire [19:0] TLB_1_xor47;
  wire [19:0] TLB_1_xor97;
  wire [19:0] TLB_1_xor98;
  wire [19:0] TLB_1_xor48;
  wire [19:0] TLB_1_xor23;
  wire [19:0] TLB_1_xor100;
  wire [19:0] TLB_1_xor49;
  wire [19:0] TLB_1_xor101;
  wire [19:0] TLB_1_xor102;
  wire [19:0] TLB_1_xor50;
  wire [19:0] TLB_1_xor24;
  wire [19:0] TLB_1_xor11;
  wire [19:0] TLB_1_xor104;
  wire [19:0] TLB_1_xor51;
  wire [19:0] TLB_1_xor105;
  wire [19:0] TLB_1_xor106;
  wire [19:0] TLB_1_xor52;
  wire [19:0] TLB_1_xor25;
  wire [19:0] TLB_1_xor107;
  wire [19:0] TLB_1_xor108;
  wire [19:0] TLB_1_xor53;
  wire [19:0] TLB_1_xor109;
  wire [19:0] TLB_1_xor110;
  wire [19:0] TLB_1_xor54;
  wire [19:0] TLB_1_xor26;
  wire [19:0] TLB_1_xor12;
  wire [19:0] TLB_1_xor5;
  wire [19:0] TLB_1_xor112;
  wire [19:0] TLB_1_xor55;
  wire [19:0] TLB_1_xor113;
  wire [19:0] TLB_1_xor114;
  wire [19:0] TLB_1_xor56;
  wire [19:0] TLB_1_xor27;
  wire [19:0] TLB_1_xor116;
  wire [19:0] TLB_1_xor57;
  wire [19:0] TLB_1_xor117;
  wire [19:0] TLB_1_xor118;
  wire [19:0] TLB_1_xor58;
  wire [19:0] TLB_1_xor28;
  wire [19:0] TLB_1_xor13;
  wire [19:0] TLB_1_xor120;
  wire [19:0] TLB_1_xor59;
  wire [19:0] TLB_1_xor121;
  wire [19:0] TLB_1_xor122;
  wire [19:0] TLB_1_xor60;
  wire [19:0] TLB_1_xor29;
  wire [19:0] TLB_1_xor123;
  wire [19:0] TLB_1_xor124;
  wire [19:0] TLB_1_xor61;
  wire [19:0] TLB_1_xor125;
  wire [19:0] TLB_1_xor126;
  wire [19:0] TLB_1_xor62;
  wire [19:0] TLB_1_xor30;
  wire [19:0] TLB_1_xor14;
  wire [19:0] TLB_1_xor6;
  wire [19:0] TLB_1_xor2;
  wire [19:0] TLB_1_xor0;
  wire [29:0] OptimizationBarrier_20_sum;
  wire [29:0] OptimizationBarrier_21_sum;
  wire [29:0] OptimizationBarrier_35_sum;
  wire [29:0] OptimizationBarrier_6_sum;
  wire [29:0] OptimizationBarrier_16_sum;
  wire [29:0] OptimizationBarrier_12_sum;
  wire [29:0] OptimizationBarrier_9_sum;
  wire [29:0] OptimizationBarrier_8_sum;
  wire [29:0] OptimizationBarrier_2_sum;
  wire [29:0] OptimizationBarrier_25_sum;
  wire [29:0] OptimizationBarrier_23_sum;
  wire [29:0] OptimizationBarrier_27_sum;
  wire [29:0] OptimizationBarrier_30_sum;
  wire [29:0] OptimizationBarrier_1_sum;
  wire [29:0] OptimizationBarrier_18_sum;
  wire [29:0] OptimizationBarrier_31_sum;
  wire [29:0] OptimizationBarrier_19_sum;
  wire [29:0] OptimizationBarrier_37_sum;
  wire [29:0] OptimizationBarrier_28_sum;
  wire [29:0] OptimizationBarrier_33_sum;
  wire [29:0] OptimizationBarrier_4_sum;
  wire [29:0] OptimizationBarrier_38_sum;
  wire [29:0] pmp_sum;
  wire [29:0] OptimizationBarrier_sum;
  wire [29:0] OptimizationBarrier_34_sum;
  wire [29:0] OptimizationBarrier_24_sum;
  wire [29:0] OptimizationBarrier_22_sum;
  wire [29:0] OptimizationBarrier_10_sum;
  wire [29:0] OptimizationBarrier_3_sum;
  wire [29:0] OptimizationBarrier_5_sum;
  wire [29:0] OptimizationBarrier_36_sum;
  wire [29:0] OptimizationBarrier_17_sum;
  wire [29:0] OptimizationBarrier_15_sum;
  wire [29:0] OptimizationBarrier_29_sum;
  wire [29:0] OptimizationBarrier_32_sum;
  wire [29:0] OptimizationBarrier_7_sum;
  wire [29:0] OptimizationBarrier_14_sum;
  wire [29:0] OptimizationBarrier_26_sum;
  wire [29:0] OptimizationBarrier_11_sum;
  wire [29:0] OptimizationBarrier_13_sum;
  wire  stopEn0;
  wire  OptimizationBarrier_34_metaAssert_wire;
  wire  OptimizationBarrier_20_metaAssert_wire;
  wire  OptimizationBarrier_6_metaAssert_wire;
  wire  OptimizationBarrier_22_metaAssert_wire;
  wire  OptimizationBarrier_14_metaAssert_wire;
  wire  OptimizationBarrier_36_metaAssert_wire;
  wire  OptimizationBarrier_37_metaAssert_wire;
  wire  OptimizationBarrier_16_metaAssert_wire;
  wire  OptimizationBarrier_35_metaAssert_wire;
  wire  OptimizationBarrier_metaAssert_wire;
  wire  OptimizationBarrier_24_metaAssert_wire;
  wire  OptimizationBarrier_32_metaAssert_wire;
  wire  pmp_metaAssert_wire;
  wire  OptimizationBarrier_33_metaAssert_wire;
  wire  OptimizationBarrier_25_metaAssert_wire;
  wire  OptimizationBarrier_4_metaAssert_wire;
  wire  OptimizationBarrier_30_metaAssert_wire;
  wire  OptimizationBarrier_23_metaAssert_wire;
  wire  OptimizationBarrier_7_metaAssert_wire;
  wire  OptimizationBarrier_10_metaAssert_wire;
  wire  OptimizationBarrier_15_metaAssert_wire;
  wire  OptimizationBarrier_8_metaAssert_wire;
  wire  OptimizationBarrier_28_metaAssert_wire;
  wire  OptimizationBarrier_3_metaAssert_wire;
  wire  OptimizationBarrier_18_metaAssert_wire;
  wire  OptimizationBarrier_2_metaAssert_wire;
  wire  OptimizationBarrier_31_metaAssert_wire;
  wire  OptimizationBarrier_26_metaAssert_wire;
  wire  OptimizationBarrier_11_metaAssert_wire;
  wire  OptimizationBarrier_19_metaAssert_wire;
  wire  OptimizationBarrier_9_metaAssert_wire;
  wire  OptimizationBarrier_1_metaAssert_wire;
  wire  OptimizationBarrier_5_metaAssert_wire;
  wire  OptimizationBarrier_12_metaAssert_wire;
  wire  OptimizationBarrier_38_metaAssert_wire;
  wire  OptimizationBarrier_17_metaAssert_wire;
  wire  OptimizationBarrier_27_metaAssert_wire;
  wire  OptimizationBarrier_29_metaAssert_wire;
  wire  OptimizationBarrier_13_metaAssert_wire;
  wire  OptimizationBarrier_21_metaAssert_wire;
  wire  TLB_1_or15;
  wire  TLB_1_or34;
  wire  TLB_1_or16;
  wire  TLB_1_or7;
  wire  TLB_1_or17;
  wire  TLB_1_or38;
  wire  TLB_1_or18;
  wire  TLB_1_or8;
  wire  TLB_1_or3;
  wire  TLB_1_or19;
  wire  TLB_1_or42;
  wire  TLB_1_or20;
  wire  TLB_1_or9;
  wire  TLB_1_or21;
  wire  TLB_1_or46;
  wire  TLB_1_or22;
  wire  TLB_1_or10;
  wire  TLB_1_or4;
  wire  TLB_1_or1;
  wire  TLB_1_or23;
  wire  TLB_1_or50;
  wire  TLB_1_or24;
  wire  TLB_1_or11;
  wire  TLB_1_or25;
  wire  TLB_1_or54;
  wire  TLB_1_or26;
  wire  TLB_1_or12;
  wire  TLB_1_or5;
  wire  TLB_1_or27;
  wire  TLB_1_or58;
  wire  TLB_1_or28;
  wire  TLB_1_or13;
  wire  TLB_1_or60;
  wire  TLB_1_or29;
  wire  TLB_1_or62;
  wire  TLB_1_or30;
  wire  TLB_1_or14;
  wire  TLB_1_or6;
  wire  TLB_1_or2;
  wire  TLB_1_or0;
  reg  TLB_1_metaAssert;
  reg [31:0] _RAND_103;
  OptimizationBarrier OptimizationBarrier ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_io_x_ppn),
    .io_x_u(OptimizationBarrier_io_x_u),
    .io_x_ae(OptimizationBarrier_io_x_ae),
    .io_x_sw(OptimizationBarrier_io_x_sw),
    .io_x_sx(OptimizationBarrier_io_x_sx),
    .io_x_sr(OptimizationBarrier_io_x_sr),
    .io_x_pw(OptimizationBarrier_io_x_pw),
    .io_x_px(OptimizationBarrier_io_x_px),
    .io_x_pr(OptimizationBarrier_io_x_pr),
    .io_x_ppp(OptimizationBarrier_io_x_ppp),
    .io_x_pal(OptimizationBarrier_io_x_pal),
    .io_x_paa(OptimizationBarrier_io_x_paa),
    .io_x_eff(OptimizationBarrier_io_x_eff),
    .io_x_c(OptimizationBarrier_io_x_c),
    .io_y_ppn(OptimizationBarrier_io_y_ppn),
    .io_y_u(OptimizationBarrier_io_y_u),
    .io_y_ae(OptimizationBarrier_io_y_ae),
    .io_y_sw(OptimizationBarrier_io_y_sw),
    .io_y_sx(OptimizationBarrier_io_y_sx),
    .io_y_sr(OptimizationBarrier_io_y_sr),
    .io_y_pw(OptimizationBarrier_io_y_pw),
    .io_y_px(OptimizationBarrier_io_y_px),
    .io_y_pr(OptimizationBarrier_io_y_pr),
    .io_y_ppp(OptimizationBarrier_io_y_ppp),
    .io_y_pal(OptimizationBarrier_io_y_pal),
    .io_y_paa(OptimizationBarrier_io_y_paa),
    .io_y_eff(OptimizationBarrier_io_y_eff),
    .io_y_c(OptimizationBarrier_io_y_c),
    .io_covSum(OptimizationBarrier_io_covSum),
    .metaAssert(OptimizationBarrier_metaAssert)
  );
  PMPChecker_2 pmp ( // @[TLB.scala 190:19]
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x),
    .io_covSum(pmp_io_covSum),
    .metaAssert(pmp_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_1 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_1_io_x_ppn),
    .io_x_u(OptimizationBarrier_1_io_x_u),
    .io_x_ae(OptimizationBarrier_1_io_x_ae),
    .io_x_sw(OptimizationBarrier_1_io_x_sw),
    .io_x_sx(OptimizationBarrier_1_io_x_sx),
    .io_x_sr(OptimizationBarrier_1_io_x_sr),
    .io_x_pw(OptimizationBarrier_1_io_x_pw),
    .io_x_px(OptimizationBarrier_1_io_x_px),
    .io_x_pr(OptimizationBarrier_1_io_x_pr),
    .io_x_ppp(OptimizationBarrier_1_io_x_ppp),
    .io_x_pal(OptimizationBarrier_1_io_x_pal),
    .io_x_paa(OptimizationBarrier_1_io_x_paa),
    .io_x_eff(OptimizationBarrier_1_io_x_eff),
    .io_x_c(OptimizationBarrier_1_io_x_c),
    .io_y_ppn(OptimizationBarrier_1_io_y_ppn),
    .io_y_u(OptimizationBarrier_1_io_y_u),
    .io_y_ae(OptimizationBarrier_1_io_y_ae),
    .io_y_sw(OptimizationBarrier_1_io_y_sw),
    .io_y_sx(OptimizationBarrier_1_io_y_sx),
    .io_y_sr(OptimizationBarrier_1_io_y_sr),
    .io_y_pw(OptimizationBarrier_1_io_y_pw),
    .io_y_px(OptimizationBarrier_1_io_y_px),
    .io_y_pr(OptimizationBarrier_1_io_y_pr),
    .io_y_ppp(OptimizationBarrier_1_io_y_ppp),
    .io_y_pal(OptimizationBarrier_1_io_y_pal),
    .io_y_paa(OptimizationBarrier_1_io_y_paa),
    .io_y_eff(OptimizationBarrier_1_io_y_eff),
    .io_y_c(OptimizationBarrier_1_io_y_c),
    .io_covSum(OptimizationBarrier_1_io_covSum),
    .metaAssert(OptimizationBarrier_1_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_2 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_2_io_x_ppn),
    .io_x_u(OptimizationBarrier_2_io_x_u),
    .io_x_ae(OptimizationBarrier_2_io_x_ae),
    .io_x_sw(OptimizationBarrier_2_io_x_sw),
    .io_x_sx(OptimizationBarrier_2_io_x_sx),
    .io_x_sr(OptimizationBarrier_2_io_x_sr),
    .io_x_pw(OptimizationBarrier_2_io_x_pw),
    .io_x_px(OptimizationBarrier_2_io_x_px),
    .io_x_pr(OptimizationBarrier_2_io_x_pr),
    .io_x_ppp(OptimizationBarrier_2_io_x_ppp),
    .io_x_pal(OptimizationBarrier_2_io_x_pal),
    .io_x_paa(OptimizationBarrier_2_io_x_paa),
    .io_x_eff(OptimizationBarrier_2_io_x_eff),
    .io_x_c(OptimizationBarrier_2_io_x_c),
    .io_y_ppn(OptimizationBarrier_2_io_y_ppn),
    .io_y_u(OptimizationBarrier_2_io_y_u),
    .io_y_ae(OptimizationBarrier_2_io_y_ae),
    .io_y_sw(OptimizationBarrier_2_io_y_sw),
    .io_y_sx(OptimizationBarrier_2_io_y_sx),
    .io_y_sr(OptimizationBarrier_2_io_y_sr),
    .io_y_pw(OptimizationBarrier_2_io_y_pw),
    .io_y_px(OptimizationBarrier_2_io_y_px),
    .io_y_pr(OptimizationBarrier_2_io_y_pr),
    .io_y_ppp(OptimizationBarrier_2_io_y_ppp),
    .io_y_pal(OptimizationBarrier_2_io_y_pal),
    .io_y_paa(OptimizationBarrier_2_io_y_paa),
    .io_y_eff(OptimizationBarrier_2_io_y_eff),
    .io_y_c(OptimizationBarrier_2_io_y_c),
    .io_covSum(OptimizationBarrier_2_io_covSum),
    .metaAssert(OptimizationBarrier_2_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_3 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_3_io_x_ppn),
    .io_x_u(OptimizationBarrier_3_io_x_u),
    .io_x_ae(OptimizationBarrier_3_io_x_ae),
    .io_x_sw(OptimizationBarrier_3_io_x_sw),
    .io_x_sx(OptimizationBarrier_3_io_x_sx),
    .io_x_sr(OptimizationBarrier_3_io_x_sr),
    .io_x_pw(OptimizationBarrier_3_io_x_pw),
    .io_x_px(OptimizationBarrier_3_io_x_px),
    .io_x_pr(OptimizationBarrier_3_io_x_pr),
    .io_x_ppp(OptimizationBarrier_3_io_x_ppp),
    .io_x_pal(OptimizationBarrier_3_io_x_pal),
    .io_x_paa(OptimizationBarrier_3_io_x_paa),
    .io_x_eff(OptimizationBarrier_3_io_x_eff),
    .io_x_c(OptimizationBarrier_3_io_x_c),
    .io_y_ppn(OptimizationBarrier_3_io_y_ppn),
    .io_y_u(OptimizationBarrier_3_io_y_u),
    .io_y_ae(OptimizationBarrier_3_io_y_ae),
    .io_y_sw(OptimizationBarrier_3_io_y_sw),
    .io_y_sx(OptimizationBarrier_3_io_y_sx),
    .io_y_sr(OptimizationBarrier_3_io_y_sr),
    .io_y_pw(OptimizationBarrier_3_io_y_pw),
    .io_y_px(OptimizationBarrier_3_io_y_px),
    .io_y_pr(OptimizationBarrier_3_io_y_pr),
    .io_y_ppp(OptimizationBarrier_3_io_y_ppp),
    .io_y_pal(OptimizationBarrier_3_io_y_pal),
    .io_y_paa(OptimizationBarrier_3_io_y_paa),
    .io_y_eff(OptimizationBarrier_3_io_y_eff),
    .io_y_c(OptimizationBarrier_3_io_y_c),
    .io_covSum(OptimizationBarrier_3_io_covSum),
    .metaAssert(OptimizationBarrier_3_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_4 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_4_io_x_ppn),
    .io_x_u(OptimizationBarrier_4_io_x_u),
    .io_x_ae(OptimizationBarrier_4_io_x_ae),
    .io_x_sw(OptimizationBarrier_4_io_x_sw),
    .io_x_sx(OptimizationBarrier_4_io_x_sx),
    .io_x_sr(OptimizationBarrier_4_io_x_sr),
    .io_x_pw(OptimizationBarrier_4_io_x_pw),
    .io_x_px(OptimizationBarrier_4_io_x_px),
    .io_x_pr(OptimizationBarrier_4_io_x_pr),
    .io_x_ppp(OptimizationBarrier_4_io_x_ppp),
    .io_x_pal(OptimizationBarrier_4_io_x_pal),
    .io_x_paa(OptimizationBarrier_4_io_x_paa),
    .io_x_eff(OptimizationBarrier_4_io_x_eff),
    .io_x_c(OptimizationBarrier_4_io_x_c),
    .io_y_ppn(OptimizationBarrier_4_io_y_ppn),
    .io_y_u(OptimizationBarrier_4_io_y_u),
    .io_y_ae(OptimizationBarrier_4_io_y_ae),
    .io_y_sw(OptimizationBarrier_4_io_y_sw),
    .io_y_sx(OptimizationBarrier_4_io_y_sx),
    .io_y_sr(OptimizationBarrier_4_io_y_sr),
    .io_y_pw(OptimizationBarrier_4_io_y_pw),
    .io_y_px(OptimizationBarrier_4_io_y_px),
    .io_y_pr(OptimizationBarrier_4_io_y_pr),
    .io_y_ppp(OptimizationBarrier_4_io_y_ppp),
    .io_y_pal(OptimizationBarrier_4_io_y_pal),
    .io_y_paa(OptimizationBarrier_4_io_y_paa),
    .io_y_eff(OptimizationBarrier_4_io_y_eff),
    .io_y_c(OptimizationBarrier_4_io_y_c),
    .io_covSum(OptimizationBarrier_4_io_covSum),
    .metaAssert(OptimizationBarrier_4_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_5 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_5_io_x_ppn),
    .io_x_u(OptimizationBarrier_5_io_x_u),
    .io_x_ae(OptimizationBarrier_5_io_x_ae),
    .io_x_sw(OptimizationBarrier_5_io_x_sw),
    .io_x_sx(OptimizationBarrier_5_io_x_sx),
    .io_x_sr(OptimizationBarrier_5_io_x_sr),
    .io_x_pw(OptimizationBarrier_5_io_x_pw),
    .io_x_px(OptimizationBarrier_5_io_x_px),
    .io_x_pr(OptimizationBarrier_5_io_x_pr),
    .io_x_ppp(OptimizationBarrier_5_io_x_ppp),
    .io_x_pal(OptimizationBarrier_5_io_x_pal),
    .io_x_paa(OptimizationBarrier_5_io_x_paa),
    .io_x_eff(OptimizationBarrier_5_io_x_eff),
    .io_x_c(OptimizationBarrier_5_io_x_c),
    .io_y_ppn(OptimizationBarrier_5_io_y_ppn),
    .io_y_u(OptimizationBarrier_5_io_y_u),
    .io_y_ae(OptimizationBarrier_5_io_y_ae),
    .io_y_sw(OptimizationBarrier_5_io_y_sw),
    .io_y_sx(OptimizationBarrier_5_io_y_sx),
    .io_y_sr(OptimizationBarrier_5_io_y_sr),
    .io_y_pw(OptimizationBarrier_5_io_y_pw),
    .io_y_px(OptimizationBarrier_5_io_y_px),
    .io_y_pr(OptimizationBarrier_5_io_y_pr),
    .io_y_ppp(OptimizationBarrier_5_io_y_ppp),
    .io_y_pal(OptimizationBarrier_5_io_y_pal),
    .io_y_paa(OptimizationBarrier_5_io_y_paa),
    .io_y_eff(OptimizationBarrier_5_io_y_eff),
    .io_y_c(OptimizationBarrier_5_io_y_c),
    .io_covSum(OptimizationBarrier_5_io_covSum),
    .metaAssert(OptimizationBarrier_5_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_6 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_6_io_x_ppn),
    .io_x_u(OptimizationBarrier_6_io_x_u),
    .io_x_ae(OptimizationBarrier_6_io_x_ae),
    .io_x_sw(OptimizationBarrier_6_io_x_sw),
    .io_x_sx(OptimizationBarrier_6_io_x_sx),
    .io_x_sr(OptimizationBarrier_6_io_x_sr),
    .io_x_pw(OptimizationBarrier_6_io_x_pw),
    .io_x_px(OptimizationBarrier_6_io_x_px),
    .io_x_pr(OptimizationBarrier_6_io_x_pr),
    .io_x_ppp(OptimizationBarrier_6_io_x_ppp),
    .io_x_pal(OptimizationBarrier_6_io_x_pal),
    .io_x_paa(OptimizationBarrier_6_io_x_paa),
    .io_x_eff(OptimizationBarrier_6_io_x_eff),
    .io_x_c(OptimizationBarrier_6_io_x_c),
    .io_y_ppn(OptimizationBarrier_6_io_y_ppn),
    .io_y_u(OptimizationBarrier_6_io_y_u),
    .io_y_ae(OptimizationBarrier_6_io_y_ae),
    .io_y_sw(OptimizationBarrier_6_io_y_sw),
    .io_y_sx(OptimizationBarrier_6_io_y_sx),
    .io_y_sr(OptimizationBarrier_6_io_y_sr),
    .io_y_pw(OptimizationBarrier_6_io_y_pw),
    .io_y_px(OptimizationBarrier_6_io_y_px),
    .io_y_pr(OptimizationBarrier_6_io_y_pr),
    .io_y_ppp(OptimizationBarrier_6_io_y_ppp),
    .io_y_pal(OptimizationBarrier_6_io_y_pal),
    .io_y_paa(OptimizationBarrier_6_io_y_paa),
    .io_y_eff(OptimizationBarrier_6_io_y_eff),
    .io_y_c(OptimizationBarrier_6_io_y_c),
    .io_covSum(OptimizationBarrier_6_io_covSum),
    .metaAssert(OptimizationBarrier_6_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_7 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_7_io_x_ppn),
    .io_x_u(OptimizationBarrier_7_io_x_u),
    .io_x_ae(OptimizationBarrier_7_io_x_ae),
    .io_x_sw(OptimizationBarrier_7_io_x_sw),
    .io_x_sx(OptimizationBarrier_7_io_x_sx),
    .io_x_sr(OptimizationBarrier_7_io_x_sr),
    .io_x_pw(OptimizationBarrier_7_io_x_pw),
    .io_x_px(OptimizationBarrier_7_io_x_px),
    .io_x_pr(OptimizationBarrier_7_io_x_pr),
    .io_x_ppp(OptimizationBarrier_7_io_x_ppp),
    .io_x_pal(OptimizationBarrier_7_io_x_pal),
    .io_x_paa(OptimizationBarrier_7_io_x_paa),
    .io_x_eff(OptimizationBarrier_7_io_x_eff),
    .io_x_c(OptimizationBarrier_7_io_x_c),
    .io_y_ppn(OptimizationBarrier_7_io_y_ppn),
    .io_y_u(OptimizationBarrier_7_io_y_u),
    .io_y_ae(OptimizationBarrier_7_io_y_ae),
    .io_y_sw(OptimizationBarrier_7_io_y_sw),
    .io_y_sx(OptimizationBarrier_7_io_y_sx),
    .io_y_sr(OptimizationBarrier_7_io_y_sr),
    .io_y_pw(OptimizationBarrier_7_io_y_pw),
    .io_y_px(OptimizationBarrier_7_io_y_px),
    .io_y_pr(OptimizationBarrier_7_io_y_pr),
    .io_y_ppp(OptimizationBarrier_7_io_y_ppp),
    .io_y_pal(OptimizationBarrier_7_io_y_pal),
    .io_y_paa(OptimizationBarrier_7_io_y_paa),
    .io_y_eff(OptimizationBarrier_7_io_y_eff),
    .io_y_c(OptimizationBarrier_7_io_y_c),
    .io_covSum(OptimizationBarrier_7_io_covSum),
    .metaAssert(OptimizationBarrier_7_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_8 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_8_io_x_ppn),
    .io_x_u(OptimizationBarrier_8_io_x_u),
    .io_x_ae(OptimizationBarrier_8_io_x_ae),
    .io_x_sw(OptimizationBarrier_8_io_x_sw),
    .io_x_sx(OptimizationBarrier_8_io_x_sx),
    .io_x_sr(OptimizationBarrier_8_io_x_sr),
    .io_x_pw(OptimizationBarrier_8_io_x_pw),
    .io_x_px(OptimizationBarrier_8_io_x_px),
    .io_x_pr(OptimizationBarrier_8_io_x_pr),
    .io_x_ppp(OptimizationBarrier_8_io_x_ppp),
    .io_x_pal(OptimizationBarrier_8_io_x_pal),
    .io_x_paa(OptimizationBarrier_8_io_x_paa),
    .io_x_eff(OptimizationBarrier_8_io_x_eff),
    .io_x_c(OptimizationBarrier_8_io_x_c),
    .io_y_ppn(OptimizationBarrier_8_io_y_ppn),
    .io_y_u(OptimizationBarrier_8_io_y_u),
    .io_y_ae(OptimizationBarrier_8_io_y_ae),
    .io_y_sw(OptimizationBarrier_8_io_y_sw),
    .io_y_sx(OptimizationBarrier_8_io_y_sx),
    .io_y_sr(OptimizationBarrier_8_io_y_sr),
    .io_y_pw(OptimizationBarrier_8_io_y_pw),
    .io_y_px(OptimizationBarrier_8_io_y_px),
    .io_y_pr(OptimizationBarrier_8_io_y_pr),
    .io_y_ppp(OptimizationBarrier_8_io_y_ppp),
    .io_y_pal(OptimizationBarrier_8_io_y_pal),
    .io_y_paa(OptimizationBarrier_8_io_y_paa),
    .io_y_eff(OptimizationBarrier_8_io_y_eff),
    .io_y_c(OptimizationBarrier_8_io_y_c),
    .io_covSum(OptimizationBarrier_8_io_covSum),
    .metaAssert(OptimizationBarrier_8_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_9 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_9_io_x_ppn),
    .io_x_u(OptimizationBarrier_9_io_x_u),
    .io_x_ae(OptimizationBarrier_9_io_x_ae),
    .io_x_sw(OptimizationBarrier_9_io_x_sw),
    .io_x_sx(OptimizationBarrier_9_io_x_sx),
    .io_x_sr(OptimizationBarrier_9_io_x_sr),
    .io_x_pw(OptimizationBarrier_9_io_x_pw),
    .io_x_px(OptimizationBarrier_9_io_x_px),
    .io_x_pr(OptimizationBarrier_9_io_x_pr),
    .io_x_ppp(OptimizationBarrier_9_io_x_ppp),
    .io_x_pal(OptimizationBarrier_9_io_x_pal),
    .io_x_paa(OptimizationBarrier_9_io_x_paa),
    .io_x_eff(OptimizationBarrier_9_io_x_eff),
    .io_x_c(OptimizationBarrier_9_io_x_c),
    .io_y_ppn(OptimizationBarrier_9_io_y_ppn),
    .io_y_u(OptimizationBarrier_9_io_y_u),
    .io_y_ae(OptimizationBarrier_9_io_y_ae),
    .io_y_sw(OptimizationBarrier_9_io_y_sw),
    .io_y_sx(OptimizationBarrier_9_io_y_sx),
    .io_y_sr(OptimizationBarrier_9_io_y_sr),
    .io_y_pw(OptimizationBarrier_9_io_y_pw),
    .io_y_px(OptimizationBarrier_9_io_y_px),
    .io_y_pr(OptimizationBarrier_9_io_y_pr),
    .io_y_ppp(OptimizationBarrier_9_io_y_ppp),
    .io_y_pal(OptimizationBarrier_9_io_y_pal),
    .io_y_paa(OptimizationBarrier_9_io_y_paa),
    .io_y_eff(OptimizationBarrier_9_io_y_eff),
    .io_y_c(OptimizationBarrier_9_io_y_c),
    .io_covSum(OptimizationBarrier_9_io_covSum),
    .metaAssert(OptimizationBarrier_9_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_10 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_10_io_x_ppn),
    .io_x_u(OptimizationBarrier_10_io_x_u),
    .io_x_ae(OptimizationBarrier_10_io_x_ae),
    .io_x_sw(OptimizationBarrier_10_io_x_sw),
    .io_x_sx(OptimizationBarrier_10_io_x_sx),
    .io_x_sr(OptimizationBarrier_10_io_x_sr),
    .io_x_pw(OptimizationBarrier_10_io_x_pw),
    .io_x_px(OptimizationBarrier_10_io_x_px),
    .io_x_pr(OptimizationBarrier_10_io_x_pr),
    .io_x_ppp(OptimizationBarrier_10_io_x_ppp),
    .io_x_pal(OptimizationBarrier_10_io_x_pal),
    .io_x_paa(OptimizationBarrier_10_io_x_paa),
    .io_x_eff(OptimizationBarrier_10_io_x_eff),
    .io_x_c(OptimizationBarrier_10_io_x_c),
    .io_y_ppn(OptimizationBarrier_10_io_y_ppn),
    .io_y_u(OptimizationBarrier_10_io_y_u),
    .io_y_ae(OptimizationBarrier_10_io_y_ae),
    .io_y_sw(OptimizationBarrier_10_io_y_sw),
    .io_y_sx(OptimizationBarrier_10_io_y_sx),
    .io_y_sr(OptimizationBarrier_10_io_y_sr),
    .io_y_pw(OptimizationBarrier_10_io_y_pw),
    .io_y_px(OptimizationBarrier_10_io_y_px),
    .io_y_pr(OptimizationBarrier_10_io_y_pr),
    .io_y_ppp(OptimizationBarrier_10_io_y_ppp),
    .io_y_pal(OptimizationBarrier_10_io_y_pal),
    .io_y_paa(OptimizationBarrier_10_io_y_paa),
    .io_y_eff(OptimizationBarrier_10_io_y_eff),
    .io_y_c(OptimizationBarrier_10_io_y_c),
    .io_covSum(OptimizationBarrier_10_io_covSum),
    .metaAssert(OptimizationBarrier_10_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_11 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_11_io_x_ppn),
    .io_x_u(OptimizationBarrier_11_io_x_u),
    .io_x_ae(OptimizationBarrier_11_io_x_ae),
    .io_x_sw(OptimizationBarrier_11_io_x_sw),
    .io_x_sx(OptimizationBarrier_11_io_x_sx),
    .io_x_sr(OptimizationBarrier_11_io_x_sr),
    .io_x_pw(OptimizationBarrier_11_io_x_pw),
    .io_x_px(OptimizationBarrier_11_io_x_px),
    .io_x_pr(OptimizationBarrier_11_io_x_pr),
    .io_x_ppp(OptimizationBarrier_11_io_x_ppp),
    .io_x_pal(OptimizationBarrier_11_io_x_pal),
    .io_x_paa(OptimizationBarrier_11_io_x_paa),
    .io_x_eff(OptimizationBarrier_11_io_x_eff),
    .io_x_c(OptimizationBarrier_11_io_x_c),
    .io_y_ppn(OptimizationBarrier_11_io_y_ppn),
    .io_y_u(OptimizationBarrier_11_io_y_u),
    .io_y_ae(OptimizationBarrier_11_io_y_ae),
    .io_y_sw(OptimizationBarrier_11_io_y_sw),
    .io_y_sx(OptimizationBarrier_11_io_y_sx),
    .io_y_sr(OptimizationBarrier_11_io_y_sr),
    .io_y_pw(OptimizationBarrier_11_io_y_pw),
    .io_y_px(OptimizationBarrier_11_io_y_px),
    .io_y_pr(OptimizationBarrier_11_io_y_pr),
    .io_y_ppp(OptimizationBarrier_11_io_y_ppp),
    .io_y_pal(OptimizationBarrier_11_io_y_pal),
    .io_y_paa(OptimizationBarrier_11_io_y_paa),
    .io_y_eff(OptimizationBarrier_11_io_y_eff),
    .io_y_c(OptimizationBarrier_11_io_y_c),
    .io_covSum(OptimizationBarrier_11_io_covSum),
    .metaAssert(OptimizationBarrier_11_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_12 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_12_io_x_ppn),
    .io_x_u(OptimizationBarrier_12_io_x_u),
    .io_x_ae(OptimizationBarrier_12_io_x_ae),
    .io_x_sw(OptimizationBarrier_12_io_x_sw),
    .io_x_sx(OptimizationBarrier_12_io_x_sx),
    .io_x_sr(OptimizationBarrier_12_io_x_sr),
    .io_x_pw(OptimizationBarrier_12_io_x_pw),
    .io_x_px(OptimizationBarrier_12_io_x_px),
    .io_x_pr(OptimizationBarrier_12_io_x_pr),
    .io_x_ppp(OptimizationBarrier_12_io_x_ppp),
    .io_x_pal(OptimizationBarrier_12_io_x_pal),
    .io_x_paa(OptimizationBarrier_12_io_x_paa),
    .io_x_eff(OptimizationBarrier_12_io_x_eff),
    .io_x_c(OptimizationBarrier_12_io_x_c),
    .io_y_ppn(OptimizationBarrier_12_io_y_ppn),
    .io_y_u(OptimizationBarrier_12_io_y_u),
    .io_y_ae(OptimizationBarrier_12_io_y_ae),
    .io_y_sw(OptimizationBarrier_12_io_y_sw),
    .io_y_sx(OptimizationBarrier_12_io_y_sx),
    .io_y_sr(OptimizationBarrier_12_io_y_sr),
    .io_y_pw(OptimizationBarrier_12_io_y_pw),
    .io_y_px(OptimizationBarrier_12_io_y_px),
    .io_y_pr(OptimizationBarrier_12_io_y_pr),
    .io_y_ppp(OptimizationBarrier_12_io_y_ppp),
    .io_y_pal(OptimizationBarrier_12_io_y_pal),
    .io_y_paa(OptimizationBarrier_12_io_y_paa),
    .io_y_eff(OptimizationBarrier_12_io_y_eff),
    .io_y_c(OptimizationBarrier_12_io_y_c),
    .io_covSum(OptimizationBarrier_12_io_covSum),
    .metaAssert(OptimizationBarrier_12_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_13 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_13_io_x_ppn),
    .io_x_u(OptimizationBarrier_13_io_x_u),
    .io_x_ae(OptimizationBarrier_13_io_x_ae),
    .io_x_sw(OptimizationBarrier_13_io_x_sw),
    .io_x_sx(OptimizationBarrier_13_io_x_sx),
    .io_x_sr(OptimizationBarrier_13_io_x_sr),
    .io_x_pw(OptimizationBarrier_13_io_x_pw),
    .io_x_px(OptimizationBarrier_13_io_x_px),
    .io_x_pr(OptimizationBarrier_13_io_x_pr),
    .io_x_ppp(OptimizationBarrier_13_io_x_ppp),
    .io_x_pal(OptimizationBarrier_13_io_x_pal),
    .io_x_paa(OptimizationBarrier_13_io_x_paa),
    .io_x_eff(OptimizationBarrier_13_io_x_eff),
    .io_x_c(OptimizationBarrier_13_io_x_c),
    .io_y_ppn(OptimizationBarrier_13_io_y_ppn),
    .io_y_u(OptimizationBarrier_13_io_y_u),
    .io_y_ae(OptimizationBarrier_13_io_y_ae),
    .io_y_sw(OptimizationBarrier_13_io_y_sw),
    .io_y_sx(OptimizationBarrier_13_io_y_sx),
    .io_y_sr(OptimizationBarrier_13_io_y_sr),
    .io_y_pw(OptimizationBarrier_13_io_y_pw),
    .io_y_px(OptimizationBarrier_13_io_y_px),
    .io_y_pr(OptimizationBarrier_13_io_y_pr),
    .io_y_ppp(OptimizationBarrier_13_io_y_ppp),
    .io_y_pal(OptimizationBarrier_13_io_y_pal),
    .io_y_paa(OptimizationBarrier_13_io_y_paa),
    .io_y_eff(OptimizationBarrier_13_io_y_eff),
    .io_y_c(OptimizationBarrier_13_io_y_c),
    .io_covSum(OptimizationBarrier_13_io_covSum),
    .metaAssert(OptimizationBarrier_13_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_14 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_14_io_x_ppn),
    .io_x_u(OptimizationBarrier_14_io_x_u),
    .io_x_ae(OptimizationBarrier_14_io_x_ae),
    .io_x_sw(OptimizationBarrier_14_io_x_sw),
    .io_x_sx(OptimizationBarrier_14_io_x_sx),
    .io_x_sr(OptimizationBarrier_14_io_x_sr),
    .io_x_pw(OptimizationBarrier_14_io_x_pw),
    .io_x_px(OptimizationBarrier_14_io_x_px),
    .io_x_pr(OptimizationBarrier_14_io_x_pr),
    .io_x_ppp(OptimizationBarrier_14_io_x_ppp),
    .io_x_pal(OptimizationBarrier_14_io_x_pal),
    .io_x_paa(OptimizationBarrier_14_io_x_paa),
    .io_x_eff(OptimizationBarrier_14_io_x_eff),
    .io_x_c(OptimizationBarrier_14_io_x_c),
    .io_y_ppn(OptimizationBarrier_14_io_y_ppn),
    .io_y_u(OptimizationBarrier_14_io_y_u),
    .io_y_ae(OptimizationBarrier_14_io_y_ae),
    .io_y_sw(OptimizationBarrier_14_io_y_sw),
    .io_y_sx(OptimizationBarrier_14_io_y_sx),
    .io_y_sr(OptimizationBarrier_14_io_y_sr),
    .io_y_pw(OptimizationBarrier_14_io_y_pw),
    .io_y_px(OptimizationBarrier_14_io_y_px),
    .io_y_pr(OptimizationBarrier_14_io_y_pr),
    .io_y_ppp(OptimizationBarrier_14_io_y_ppp),
    .io_y_pal(OptimizationBarrier_14_io_y_pal),
    .io_y_paa(OptimizationBarrier_14_io_y_paa),
    .io_y_eff(OptimizationBarrier_14_io_y_eff),
    .io_y_c(OptimizationBarrier_14_io_y_c),
    .io_covSum(OptimizationBarrier_14_io_covSum),
    .metaAssert(OptimizationBarrier_14_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_15 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_15_io_x_ppn),
    .io_x_u(OptimizationBarrier_15_io_x_u),
    .io_x_ae(OptimizationBarrier_15_io_x_ae),
    .io_x_sw(OptimizationBarrier_15_io_x_sw),
    .io_x_sx(OptimizationBarrier_15_io_x_sx),
    .io_x_sr(OptimizationBarrier_15_io_x_sr),
    .io_x_pw(OptimizationBarrier_15_io_x_pw),
    .io_x_px(OptimizationBarrier_15_io_x_px),
    .io_x_pr(OptimizationBarrier_15_io_x_pr),
    .io_x_ppp(OptimizationBarrier_15_io_x_ppp),
    .io_x_pal(OptimizationBarrier_15_io_x_pal),
    .io_x_paa(OptimizationBarrier_15_io_x_paa),
    .io_x_eff(OptimizationBarrier_15_io_x_eff),
    .io_x_c(OptimizationBarrier_15_io_x_c),
    .io_y_ppn(OptimizationBarrier_15_io_y_ppn),
    .io_y_u(OptimizationBarrier_15_io_y_u),
    .io_y_ae(OptimizationBarrier_15_io_y_ae),
    .io_y_sw(OptimizationBarrier_15_io_y_sw),
    .io_y_sx(OptimizationBarrier_15_io_y_sx),
    .io_y_sr(OptimizationBarrier_15_io_y_sr),
    .io_y_pw(OptimizationBarrier_15_io_y_pw),
    .io_y_px(OptimizationBarrier_15_io_y_px),
    .io_y_pr(OptimizationBarrier_15_io_y_pr),
    .io_y_ppp(OptimizationBarrier_15_io_y_ppp),
    .io_y_pal(OptimizationBarrier_15_io_y_pal),
    .io_y_paa(OptimizationBarrier_15_io_y_paa),
    .io_y_eff(OptimizationBarrier_15_io_y_eff),
    .io_y_c(OptimizationBarrier_15_io_y_c),
    .io_covSum(OptimizationBarrier_15_io_covSum),
    .metaAssert(OptimizationBarrier_15_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_16 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_16_io_x_ppn),
    .io_x_u(OptimizationBarrier_16_io_x_u),
    .io_x_ae(OptimizationBarrier_16_io_x_ae),
    .io_x_sw(OptimizationBarrier_16_io_x_sw),
    .io_x_sx(OptimizationBarrier_16_io_x_sx),
    .io_x_sr(OptimizationBarrier_16_io_x_sr),
    .io_x_pw(OptimizationBarrier_16_io_x_pw),
    .io_x_px(OptimizationBarrier_16_io_x_px),
    .io_x_pr(OptimizationBarrier_16_io_x_pr),
    .io_x_ppp(OptimizationBarrier_16_io_x_ppp),
    .io_x_pal(OptimizationBarrier_16_io_x_pal),
    .io_x_paa(OptimizationBarrier_16_io_x_paa),
    .io_x_eff(OptimizationBarrier_16_io_x_eff),
    .io_x_c(OptimizationBarrier_16_io_x_c),
    .io_y_ppn(OptimizationBarrier_16_io_y_ppn),
    .io_y_u(OptimizationBarrier_16_io_y_u),
    .io_y_ae(OptimizationBarrier_16_io_y_ae),
    .io_y_sw(OptimizationBarrier_16_io_y_sw),
    .io_y_sx(OptimizationBarrier_16_io_y_sx),
    .io_y_sr(OptimizationBarrier_16_io_y_sr),
    .io_y_pw(OptimizationBarrier_16_io_y_pw),
    .io_y_px(OptimizationBarrier_16_io_y_px),
    .io_y_pr(OptimizationBarrier_16_io_y_pr),
    .io_y_ppp(OptimizationBarrier_16_io_y_ppp),
    .io_y_pal(OptimizationBarrier_16_io_y_pal),
    .io_y_paa(OptimizationBarrier_16_io_y_paa),
    .io_y_eff(OptimizationBarrier_16_io_y_eff),
    .io_y_c(OptimizationBarrier_16_io_y_c),
    .io_covSum(OptimizationBarrier_16_io_covSum),
    .metaAssert(OptimizationBarrier_16_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_17 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_17_io_x_ppn),
    .io_x_u(OptimizationBarrier_17_io_x_u),
    .io_x_ae(OptimizationBarrier_17_io_x_ae),
    .io_x_sw(OptimizationBarrier_17_io_x_sw),
    .io_x_sx(OptimizationBarrier_17_io_x_sx),
    .io_x_sr(OptimizationBarrier_17_io_x_sr),
    .io_x_pw(OptimizationBarrier_17_io_x_pw),
    .io_x_px(OptimizationBarrier_17_io_x_px),
    .io_x_pr(OptimizationBarrier_17_io_x_pr),
    .io_x_ppp(OptimizationBarrier_17_io_x_ppp),
    .io_x_pal(OptimizationBarrier_17_io_x_pal),
    .io_x_paa(OptimizationBarrier_17_io_x_paa),
    .io_x_eff(OptimizationBarrier_17_io_x_eff),
    .io_x_c(OptimizationBarrier_17_io_x_c),
    .io_y_ppn(OptimizationBarrier_17_io_y_ppn),
    .io_y_u(OptimizationBarrier_17_io_y_u),
    .io_y_ae(OptimizationBarrier_17_io_y_ae),
    .io_y_sw(OptimizationBarrier_17_io_y_sw),
    .io_y_sx(OptimizationBarrier_17_io_y_sx),
    .io_y_sr(OptimizationBarrier_17_io_y_sr),
    .io_y_pw(OptimizationBarrier_17_io_y_pw),
    .io_y_px(OptimizationBarrier_17_io_y_px),
    .io_y_pr(OptimizationBarrier_17_io_y_pr),
    .io_y_ppp(OptimizationBarrier_17_io_y_ppp),
    .io_y_pal(OptimizationBarrier_17_io_y_pal),
    .io_y_paa(OptimizationBarrier_17_io_y_paa),
    .io_y_eff(OptimizationBarrier_17_io_y_eff),
    .io_y_c(OptimizationBarrier_17_io_y_c),
    .io_covSum(OptimizationBarrier_17_io_covSum),
    .metaAssert(OptimizationBarrier_17_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_18 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_18_io_x_ppn),
    .io_x_u(OptimizationBarrier_18_io_x_u),
    .io_x_ae(OptimizationBarrier_18_io_x_ae),
    .io_x_sw(OptimizationBarrier_18_io_x_sw),
    .io_x_sx(OptimizationBarrier_18_io_x_sx),
    .io_x_sr(OptimizationBarrier_18_io_x_sr),
    .io_x_pw(OptimizationBarrier_18_io_x_pw),
    .io_x_px(OptimizationBarrier_18_io_x_px),
    .io_x_pr(OptimizationBarrier_18_io_x_pr),
    .io_x_ppp(OptimizationBarrier_18_io_x_ppp),
    .io_x_pal(OptimizationBarrier_18_io_x_pal),
    .io_x_paa(OptimizationBarrier_18_io_x_paa),
    .io_x_eff(OptimizationBarrier_18_io_x_eff),
    .io_x_c(OptimizationBarrier_18_io_x_c),
    .io_y_ppn(OptimizationBarrier_18_io_y_ppn),
    .io_y_u(OptimizationBarrier_18_io_y_u),
    .io_y_ae(OptimizationBarrier_18_io_y_ae),
    .io_y_sw(OptimizationBarrier_18_io_y_sw),
    .io_y_sx(OptimizationBarrier_18_io_y_sx),
    .io_y_sr(OptimizationBarrier_18_io_y_sr),
    .io_y_pw(OptimizationBarrier_18_io_y_pw),
    .io_y_px(OptimizationBarrier_18_io_y_px),
    .io_y_pr(OptimizationBarrier_18_io_y_pr),
    .io_y_ppp(OptimizationBarrier_18_io_y_ppp),
    .io_y_pal(OptimizationBarrier_18_io_y_pal),
    .io_y_paa(OptimizationBarrier_18_io_y_paa),
    .io_y_eff(OptimizationBarrier_18_io_y_eff),
    .io_y_c(OptimizationBarrier_18_io_y_c),
    .io_covSum(OptimizationBarrier_18_io_covSum),
    .metaAssert(OptimizationBarrier_18_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_19 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_19_io_x_ppn),
    .io_x_u(OptimizationBarrier_19_io_x_u),
    .io_x_ae(OptimizationBarrier_19_io_x_ae),
    .io_x_sw(OptimizationBarrier_19_io_x_sw),
    .io_x_sx(OptimizationBarrier_19_io_x_sx),
    .io_x_sr(OptimizationBarrier_19_io_x_sr),
    .io_x_pw(OptimizationBarrier_19_io_x_pw),
    .io_x_px(OptimizationBarrier_19_io_x_px),
    .io_x_pr(OptimizationBarrier_19_io_x_pr),
    .io_x_ppp(OptimizationBarrier_19_io_x_ppp),
    .io_x_pal(OptimizationBarrier_19_io_x_pal),
    .io_x_paa(OptimizationBarrier_19_io_x_paa),
    .io_x_eff(OptimizationBarrier_19_io_x_eff),
    .io_x_c(OptimizationBarrier_19_io_x_c),
    .io_y_ppn(OptimizationBarrier_19_io_y_ppn),
    .io_y_u(OptimizationBarrier_19_io_y_u),
    .io_y_ae(OptimizationBarrier_19_io_y_ae),
    .io_y_sw(OptimizationBarrier_19_io_y_sw),
    .io_y_sx(OptimizationBarrier_19_io_y_sx),
    .io_y_sr(OptimizationBarrier_19_io_y_sr),
    .io_y_pw(OptimizationBarrier_19_io_y_pw),
    .io_y_px(OptimizationBarrier_19_io_y_px),
    .io_y_pr(OptimizationBarrier_19_io_y_pr),
    .io_y_ppp(OptimizationBarrier_19_io_y_ppp),
    .io_y_pal(OptimizationBarrier_19_io_y_pal),
    .io_y_paa(OptimizationBarrier_19_io_y_paa),
    .io_y_eff(OptimizationBarrier_19_io_y_eff),
    .io_y_c(OptimizationBarrier_19_io_y_c),
    .io_covSum(OptimizationBarrier_19_io_covSum),
    .metaAssert(OptimizationBarrier_19_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_20 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_20_io_x_ppn),
    .io_x_u(OptimizationBarrier_20_io_x_u),
    .io_x_ae(OptimizationBarrier_20_io_x_ae),
    .io_x_sw(OptimizationBarrier_20_io_x_sw),
    .io_x_sx(OptimizationBarrier_20_io_x_sx),
    .io_x_sr(OptimizationBarrier_20_io_x_sr),
    .io_x_pw(OptimizationBarrier_20_io_x_pw),
    .io_x_px(OptimizationBarrier_20_io_x_px),
    .io_x_pr(OptimizationBarrier_20_io_x_pr),
    .io_x_ppp(OptimizationBarrier_20_io_x_ppp),
    .io_x_pal(OptimizationBarrier_20_io_x_pal),
    .io_x_paa(OptimizationBarrier_20_io_x_paa),
    .io_x_eff(OptimizationBarrier_20_io_x_eff),
    .io_x_c(OptimizationBarrier_20_io_x_c),
    .io_y_ppn(OptimizationBarrier_20_io_y_ppn),
    .io_y_u(OptimizationBarrier_20_io_y_u),
    .io_y_ae(OptimizationBarrier_20_io_y_ae),
    .io_y_sw(OptimizationBarrier_20_io_y_sw),
    .io_y_sx(OptimizationBarrier_20_io_y_sx),
    .io_y_sr(OptimizationBarrier_20_io_y_sr),
    .io_y_pw(OptimizationBarrier_20_io_y_pw),
    .io_y_px(OptimizationBarrier_20_io_y_px),
    .io_y_pr(OptimizationBarrier_20_io_y_pr),
    .io_y_ppp(OptimizationBarrier_20_io_y_ppp),
    .io_y_pal(OptimizationBarrier_20_io_y_pal),
    .io_y_paa(OptimizationBarrier_20_io_y_paa),
    .io_y_eff(OptimizationBarrier_20_io_y_eff),
    .io_y_c(OptimizationBarrier_20_io_y_c),
    .io_covSum(OptimizationBarrier_20_io_covSum),
    .metaAssert(OptimizationBarrier_20_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_21 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_21_io_x_ppn),
    .io_x_u(OptimizationBarrier_21_io_x_u),
    .io_x_ae(OptimizationBarrier_21_io_x_ae),
    .io_x_sw(OptimizationBarrier_21_io_x_sw),
    .io_x_sx(OptimizationBarrier_21_io_x_sx),
    .io_x_sr(OptimizationBarrier_21_io_x_sr),
    .io_x_pw(OptimizationBarrier_21_io_x_pw),
    .io_x_px(OptimizationBarrier_21_io_x_px),
    .io_x_pr(OptimizationBarrier_21_io_x_pr),
    .io_x_ppp(OptimizationBarrier_21_io_x_ppp),
    .io_x_pal(OptimizationBarrier_21_io_x_pal),
    .io_x_paa(OptimizationBarrier_21_io_x_paa),
    .io_x_eff(OptimizationBarrier_21_io_x_eff),
    .io_x_c(OptimizationBarrier_21_io_x_c),
    .io_y_ppn(OptimizationBarrier_21_io_y_ppn),
    .io_y_u(OptimizationBarrier_21_io_y_u),
    .io_y_ae(OptimizationBarrier_21_io_y_ae),
    .io_y_sw(OptimizationBarrier_21_io_y_sw),
    .io_y_sx(OptimizationBarrier_21_io_y_sx),
    .io_y_sr(OptimizationBarrier_21_io_y_sr),
    .io_y_pw(OptimizationBarrier_21_io_y_pw),
    .io_y_px(OptimizationBarrier_21_io_y_px),
    .io_y_pr(OptimizationBarrier_21_io_y_pr),
    .io_y_ppp(OptimizationBarrier_21_io_y_ppp),
    .io_y_pal(OptimizationBarrier_21_io_y_pal),
    .io_y_paa(OptimizationBarrier_21_io_y_paa),
    .io_y_eff(OptimizationBarrier_21_io_y_eff),
    .io_y_c(OptimizationBarrier_21_io_y_c),
    .io_covSum(OptimizationBarrier_21_io_covSum),
    .metaAssert(OptimizationBarrier_21_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_22 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_22_io_x_ppn),
    .io_x_u(OptimizationBarrier_22_io_x_u),
    .io_x_ae(OptimizationBarrier_22_io_x_ae),
    .io_x_sw(OptimizationBarrier_22_io_x_sw),
    .io_x_sx(OptimizationBarrier_22_io_x_sx),
    .io_x_sr(OptimizationBarrier_22_io_x_sr),
    .io_x_pw(OptimizationBarrier_22_io_x_pw),
    .io_x_px(OptimizationBarrier_22_io_x_px),
    .io_x_pr(OptimizationBarrier_22_io_x_pr),
    .io_x_ppp(OptimizationBarrier_22_io_x_ppp),
    .io_x_pal(OptimizationBarrier_22_io_x_pal),
    .io_x_paa(OptimizationBarrier_22_io_x_paa),
    .io_x_eff(OptimizationBarrier_22_io_x_eff),
    .io_x_c(OptimizationBarrier_22_io_x_c),
    .io_y_ppn(OptimizationBarrier_22_io_y_ppn),
    .io_y_u(OptimizationBarrier_22_io_y_u),
    .io_y_ae(OptimizationBarrier_22_io_y_ae),
    .io_y_sw(OptimizationBarrier_22_io_y_sw),
    .io_y_sx(OptimizationBarrier_22_io_y_sx),
    .io_y_sr(OptimizationBarrier_22_io_y_sr),
    .io_y_pw(OptimizationBarrier_22_io_y_pw),
    .io_y_px(OptimizationBarrier_22_io_y_px),
    .io_y_pr(OptimizationBarrier_22_io_y_pr),
    .io_y_ppp(OptimizationBarrier_22_io_y_ppp),
    .io_y_pal(OptimizationBarrier_22_io_y_pal),
    .io_y_paa(OptimizationBarrier_22_io_y_paa),
    .io_y_eff(OptimizationBarrier_22_io_y_eff),
    .io_y_c(OptimizationBarrier_22_io_y_c),
    .io_covSum(OptimizationBarrier_22_io_covSum),
    .metaAssert(OptimizationBarrier_22_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_23 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_23_io_x_ppn),
    .io_x_u(OptimizationBarrier_23_io_x_u),
    .io_x_ae(OptimizationBarrier_23_io_x_ae),
    .io_x_sw(OptimizationBarrier_23_io_x_sw),
    .io_x_sx(OptimizationBarrier_23_io_x_sx),
    .io_x_sr(OptimizationBarrier_23_io_x_sr),
    .io_x_pw(OptimizationBarrier_23_io_x_pw),
    .io_x_px(OptimizationBarrier_23_io_x_px),
    .io_x_pr(OptimizationBarrier_23_io_x_pr),
    .io_x_ppp(OptimizationBarrier_23_io_x_ppp),
    .io_x_pal(OptimizationBarrier_23_io_x_pal),
    .io_x_paa(OptimizationBarrier_23_io_x_paa),
    .io_x_eff(OptimizationBarrier_23_io_x_eff),
    .io_x_c(OptimizationBarrier_23_io_x_c),
    .io_y_ppn(OptimizationBarrier_23_io_y_ppn),
    .io_y_u(OptimizationBarrier_23_io_y_u),
    .io_y_ae(OptimizationBarrier_23_io_y_ae),
    .io_y_sw(OptimizationBarrier_23_io_y_sw),
    .io_y_sx(OptimizationBarrier_23_io_y_sx),
    .io_y_sr(OptimizationBarrier_23_io_y_sr),
    .io_y_pw(OptimizationBarrier_23_io_y_pw),
    .io_y_px(OptimizationBarrier_23_io_y_px),
    .io_y_pr(OptimizationBarrier_23_io_y_pr),
    .io_y_ppp(OptimizationBarrier_23_io_y_ppp),
    .io_y_pal(OptimizationBarrier_23_io_y_pal),
    .io_y_paa(OptimizationBarrier_23_io_y_paa),
    .io_y_eff(OptimizationBarrier_23_io_y_eff),
    .io_y_c(OptimizationBarrier_23_io_y_c),
    .io_covSum(OptimizationBarrier_23_io_covSum),
    .metaAssert(OptimizationBarrier_23_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_24 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_24_io_x_ppn),
    .io_x_u(OptimizationBarrier_24_io_x_u),
    .io_x_ae(OptimizationBarrier_24_io_x_ae),
    .io_x_sw(OptimizationBarrier_24_io_x_sw),
    .io_x_sx(OptimizationBarrier_24_io_x_sx),
    .io_x_sr(OptimizationBarrier_24_io_x_sr),
    .io_x_pw(OptimizationBarrier_24_io_x_pw),
    .io_x_px(OptimizationBarrier_24_io_x_px),
    .io_x_pr(OptimizationBarrier_24_io_x_pr),
    .io_x_ppp(OptimizationBarrier_24_io_x_ppp),
    .io_x_pal(OptimizationBarrier_24_io_x_pal),
    .io_x_paa(OptimizationBarrier_24_io_x_paa),
    .io_x_eff(OptimizationBarrier_24_io_x_eff),
    .io_x_c(OptimizationBarrier_24_io_x_c),
    .io_y_ppn(OptimizationBarrier_24_io_y_ppn),
    .io_y_u(OptimizationBarrier_24_io_y_u),
    .io_y_ae(OptimizationBarrier_24_io_y_ae),
    .io_y_sw(OptimizationBarrier_24_io_y_sw),
    .io_y_sx(OptimizationBarrier_24_io_y_sx),
    .io_y_sr(OptimizationBarrier_24_io_y_sr),
    .io_y_pw(OptimizationBarrier_24_io_y_pw),
    .io_y_px(OptimizationBarrier_24_io_y_px),
    .io_y_pr(OptimizationBarrier_24_io_y_pr),
    .io_y_ppp(OptimizationBarrier_24_io_y_ppp),
    .io_y_pal(OptimizationBarrier_24_io_y_pal),
    .io_y_paa(OptimizationBarrier_24_io_y_paa),
    .io_y_eff(OptimizationBarrier_24_io_y_eff),
    .io_y_c(OptimizationBarrier_24_io_y_c),
    .io_covSum(OptimizationBarrier_24_io_covSum),
    .metaAssert(OptimizationBarrier_24_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_25 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_25_io_x_ppn),
    .io_x_u(OptimizationBarrier_25_io_x_u),
    .io_x_ae(OptimizationBarrier_25_io_x_ae),
    .io_x_sw(OptimizationBarrier_25_io_x_sw),
    .io_x_sx(OptimizationBarrier_25_io_x_sx),
    .io_x_sr(OptimizationBarrier_25_io_x_sr),
    .io_x_pw(OptimizationBarrier_25_io_x_pw),
    .io_x_px(OptimizationBarrier_25_io_x_px),
    .io_x_pr(OptimizationBarrier_25_io_x_pr),
    .io_x_ppp(OptimizationBarrier_25_io_x_ppp),
    .io_x_pal(OptimizationBarrier_25_io_x_pal),
    .io_x_paa(OptimizationBarrier_25_io_x_paa),
    .io_x_eff(OptimizationBarrier_25_io_x_eff),
    .io_x_c(OptimizationBarrier_25_io_x_c),
    .io_y_ppn(OptimizationBarrier_25_io_y_ppn),
    .io_y_u(OptimizationBarrier_25_io_y_u),
    .io_y_ae(OptimizationBarrier_25_io_y_ae),
    .io_y_sw(OptimizationBarrier_25_io_y_sw),
    .io_y_sx(OptimizationBarrier_25_io_y_sx),
    .io_y_sr(OptimizationBarrier_25_io_y_sr),
    .io_y_pw(OptimizationBarrier_25_io_y_pw),
    .io_y_px(OptimizationBarrier_25_io_y_px),
    .io_y_pr(OptimizationBarrier_25_io_y_pr),
    .io_y_ppp(OptimizationBarrier_25_io_y_ppp),
    .io_y_pal(OptimizationBarrier_25_io_y_pal),
    .io_y_paa(OptimizationBarrier_25_io_y_paa),
    .io_y_eff(OptimizationBarrier_25_io_y_eff),
    .io_y_c(OptimizationBarrier_25_io_y_c),
    .io_covSum(OptimizationBarrier_25_io_covSum),
    .metaAssert(OptimizationBarrier_25_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_26 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_26_io_x_ppn),
    .io_x_u(OptimizationBarrier_26_io_x_u),
    .io_x_ae(OptimizationBarrier_26_io_x_ae),
    .io_x_sw(OptimizationBarrier_26_io_x_sw),
    .io_x_sx(OptimizationBarrier_26_io_x_sx),
    .io_x_sr(OptimizationBarrier_26_io_x_sr),
    .io_x_pw(OptimizationBarrier_26_io_x_pw),
    .io_x_px(OptimizationBarrier_26_io_x_px),
    .io_x_pr(OptimizationBarrier_26_io_x_pr),
    .io_x_ppp(OptimizationBarrier_26_io_x_ppp),
    .io_x_pal(OptimizationBarrier_26_io_x_pal),
    .io_x_paa(OptimizationBarrier_26_io_x_paa),
    .io_x_eff(OptimizationBarrier_26_io_x_eff),
    .io_x_c(OptimizationBarrier_26_io_x_c),
    .io_y_ppn(OptimizationBarrier_26_io_y_ppn),
    .io_y_u(OptimizationBarrier_26_io_y_u),
    .io_y_ae(OptimizationBarrier_26_io_y_ae),
    .io_y_sw(OptimizationBarrier_26_io_y_sw),
    .io_y_sx(OptimizationBarrier_26_io_y_sx),
    .io_y_sr(OptimizationBarrier_26_io_y_sr),
    .io_y_pw(OptimizationBarrier_26_io_y_pw),
    .io_y_px(OptimizationBarrier_26_io_y_px),
    .io_y_pr(OptimizationBarrier_26_io_y_pr),
    .io_y_ppp(OptimizationBarrier_26_io_y_ppp),
    .io_y_pal(OptimizationBarrier_26_io_y_pal),
    .io_y_paa(OptimizationBarrier_26_io_y_paa),
    .io_y_eff(OptimizationBarrier_26_io_y_eff),
    .io_y_c(OptimizationBarrier_26_io_y_c),
    .io_covSum(OptimizationBarrier_26_io_covSum),
    .metaAssert(OptimizationBarrier_26_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_27 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_27_io_x_ppn),
    .io_x_u(OptimizationBarrier_27_io_x_u),
    .io_x_ae(OptimizationBarrier_27_io_x_ae),
    .io_x_sw(OptimizationBarrier_27_io_x_sw),
    .io_x_sx(OptimizationBarrier_27_io_x_sx),
    .io_x_sr(OptimizationBarrier_27_io_x_sr),
    .io_x_pw(OptimizationBarrier_27_io_x_pw),
    .io_x_px(OptimizationBarrier_27_io_x_px),
    .io_x_pr(OptimizationBarrier_27_io_x_pr),
    .io_x_ppp(OptimizationBarrier_27_io_x_ppp),
    .io_x_pal(OptimizationBarrier_27_io_x_pal),
    .io_x_paa(OptimizationBarrier_27_io_x_paa),
    .io_x_eff(OptimizationBarrier_27_io_x_eff),
    .io_x_c(OptimizationBarrier_27_io_x_c),
    .io_y_ppn(OptimizationBarrier_27_io_y_ppn),
    .io_y_u(OptimizationBarrier_27_io_y_u),
    .io_y_ae(OptimizationBarrier_27_io_y_ae),
    .io_y_sw(OptimizationBarrier_27_io_y_sw),
    .io_y_sx(OptimizationBarrier_27_io_y_sx),
    .io_y_sr(OptimizationBarrier_27_io_y_sr),
    .io_y_pw(OptimizationBarrier_27_io_y_pw),
    .io_y_px(OptimizationBarrier_27_io_y_px),
    .io_y_pr(OptimizationBarrier_27_io_y_pr),
    .io_y_ppp(OptimizationBarrier_27_io_y_ppp),
    .io_y_pal(OptimizationBarrier_27_io_y_pal),
    .io_y_paa(OptimizationBarrier_27_io_y_paa),
    .io_y_eff(OptimizationBarrier_27_io_y_eff),
    .io_y_c(OptimizationBarrier_27_io_y_c),
    .io_covSum(OptimizationBarrier_27_io_covSum),
    .metaAssert(OptimizationBarrier_27_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_28 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_28_io_x_ppn),
    .io_x_u(OptimizationBarrier_28_io_x_u),
    .io_x_ae(OptimizationBarrier_28_io_x_ae),
    .io_x_sw(OptimizationBarrier_28_io_x_sw),
    .io_x_sx(OptimizationBarrier_28_io_x_sx),
    .io_x_sr(OptimizationBarrier_28_io_x_sr),
    .io_x_pw(OptimizationBarrier_28_io_x_pw),
    .io_x_px(OptimizationBarrier_28_io_x_px),
    .io_x_pr(OptimizationBarrier_28_io_x_pr),
    .io_x_ppp(OptimizationBarrier_28_io_x_ppp),
    .io_x_pal(OptimizationBarrier_28_io_x_pal),
    .io_x_paa(OptimizationBarrier_28_io_x_paa),
    .io_x_eff(OptimizationBarrier_28_io_x_eff),
    .io_x_c(OptimizationBarrier_28_io_x_c),
    .io_y_ppn(OptimizationBarrier_28_io_y_ppn),
    .io_y_u(OptimizationBarrier_28_io_y_u),
    .io_y_ae(OptimizationBarrier_28_io_y_ae),
    .io_y_sw(OptimizationBarrier_28_io_y_sw),
    .io_y_sx(OptimizationBarrier_28_io_y_sx),
    .io_y_sr(OptimizationBarrier_28_io_y_sr),
    .io_y_pw(OptimizationBarrier_28_io_y_pw),
    .io_y_px(OptimizationBarrier_28_io_y_px),
    .io_y_pr(OptimizationBarrier_28_io_y_pr),
    .io_y_ppp(OptimizationBarrier_28_io_y_ppp),
    .io_y_pal(OptimizationBarrier_28_io_y_pal),
    .io_y_paa(OptimizationBarrier_28_io_y_paa),
    .io_y_eff(OptimizationBarrier_28_io_y_eff),
    .io_y_c(OptimizationBarrier_28_io_y_c),
    .io_covSum(OptimizationBarrier_28_io_covSum),
    .metaAssert(OptimizationBarrier_28_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_29 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_29_io_x_ppn),
    .io_x_u(OptimizationBarrier_29_io_x_u),
    .io_x_ae(OptimizationBarrier_29_io_x_ae),
    .io_x_sw(OptimizationBarrier_29_io_x_sw),
    .io_x_sx(OptimizationBarrier_29_io_x_sx),
    .io_x_sr(OptimizationBarrier_29_io_x_sr),
    .io_x_pw(OptimizationBarrier_29_io_x_pw),
    .io_x_px(OptimizationBarrier_29_io_x_px),
    .io_x_pr(OptimizationBarrier_29_io_x_pr),
    .io_x_ppp(OptimizationBarrier_29_io_x_ppp),
    .io_x_pal(OptimizationBarrier_29_io_x_pal),
    .io_x_paa(OptimizationBarrier_29_io_x_paa),
    .io_x_eff(OptimizationBarrier_29_io_x_eff),
    .io_x_c(OptimizationBarrier_29_io_x_c),
    .io_y_ppn(OptimizationBarrier_29_io_y_ppn),
    .io_y_u(OptimizationBarrier_29_io_y_u),
    .io_y_ae(OptimizationBarrier_29_io_y_ae),
    .io_y_sw(OptimizationBarrier_29_io_y_sw),
    .io_y_sx(OptimizationBarrier_29_io_y_sx),
    .io_y_sr(OptimizationBarrier_29_io_y_sr),
    .io_y_pw(OptimizationBarrier_29_io_y_pw),
    .io_y_px(OptimizationBarrier_29_io_y_px),
    .io_y_pr(OptimizationBarrier_29_io_y_pr),
    .io_y_ppp(OptimizationBarrier_29_io_y_ppp),
    .io_y_pal(OptimizationBarrier_29_io_y_pal),
    .io_y_paa(OptimizationBarrier_29_io_y_paa),
    .io_y_eff(OptimizationBarrier_29_io_y_eff),
    .io_y_c(OptimizationBarrier_29_io_y_c),
    .io_covSum(OptimizationBarrier_29_io_covSum),
    .metaAssert(OptimizationBarrier_29_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_30 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_30_io_x_ppn),
    .io_x_u(OptimizationBarrier_30_io_x_u),
    .io_x_ae(OptimizationBarrier_30_io_x_ae),
    .io_x_sw(OptimizationBarrier_30_io_x_sw),
    .io_x_sx(OptimizationBarrier_30_io_x_sx),
    .io_x_sr(OptimizationBarrier_30_io_x_sr),
    .io_x_pw(OptimizationBarrier_30_io_x_pw),
    .io_x_px(OptimizationBarrier_30_io_x_px),
    .io_x_pr(OptimizationBarrier_30_io_x_pr),
    .io_x_ppp(OptimizationBarrier_30_io_x_ppp),
    .io_x_pal(OptimizationBarrier_30_io_x_pal),
    .io_x_paa(OptimizationBarrier_30_io_x_paa),
    .io_x_eff(OptimizationBarrier_30_io_x_eff),
    .io_x_c(OptimizationBarrier_30_io_x_c),
    .io_y_ppn(OptimizationBarrier_30_io_y_ppn),
    .io_y_u(OptimizationBarrier_30_io_y_u),
    .io_y_ae(OptimizationBarrier_30_io_y_ae),
    .io_y_sw(OptimizationBarrier_30_io_y_sw),
    .io_y_sx(OptimizationBarrier_30_io_y_sx),
    .io_y_sr(OptimizationBarrier_30_io_y_sr),
    .io_y_pw(OptimizationBarrier_30_io_y_pw),
    .io_y_px(OptimizationBarrier_30_io_y_px),
    .io_y_pr(OptimizationBarrier_30_io_y_pr),
    .io_y_ppp(OptimizationBarrier_30_io_y_ppp),
    .io_y_pal(OptimizationBarrier_30_io_y_pal),
    .io_y_paa(OptimizationBarrier_30_io_y_paa),
    .io_y_eff(OptimizationBarrier_30_io_y_eff),
    .io_y_c(OptimizationBarrier_30_io_y_c),
    .io_covSum(OptimizationBarrier_30_io_covSum),
    .metaAssert(OptimizationBarrier_30_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_31 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_31_io_x_ppn),
    .io_x_u(OptimizationBarrier_31_io_x_u),
    .io_x_ae(OptimizationBarrier_31_io_x_ae),
    .io_x_sw(OptimizationBarrier_31_io_x_sw),
    .io_x_sx(OptimizationBarrier_31_io_x_sx),
    .io_x_sr(OptimizationBarrier_31_io_x_sr),
    .io_x_pw(OptimizationBarrier_31_io_x_pw),
    .io_x_px(OptimizationBarrier_31_io_x_px),
    .io_x_pr(OptimizationBarrier_31_io_x_pr),
    .io_x_ppp(OptimizationBarrier_31_io_x_ppp),
    .io_x_pal(OptimizationBarrier_31_io_x_pal),
    .io_x_paa(OptimizationBarrier_31_io_x_paa),
    .io_x_eff(OptimizationBarrier_31_io_x_eff),
    .io_x_c(OptimizationBarrier_31_io_x_c),
    .io_y_ppn(OptimizationBarrier_31_io_y_ppn),
    .io_y_u(OptimizationBarrier_31_io_y_u),
    .io_y_ae(OptimizationBarrier_31_io_y_ae),
    .io_y_sw(OptimizationBarrier_31_io_y_sw),
    .io_y_sx(OptimizationBarrier_31_io_y_sx),
    .io_y_sr(OptimizationBarrier_31_io_y_sr),
    .io_y_pw(OptimizationBarrier_31_io_y_pw),
    .io_y_px(OptimizationBarrier_31_io_y_px),
    .io_y_pr(OptimizationBarrier_31_io_y_pr),
    .io_y_ppp(OptimizationBarrier_31_io_y_ppp),
    .io_y_pal(OptimizationBarrier_31_io_y_pal),
    .io_y_paa(OptimizationBarrier_31_io_y_paa),
    .io_y_eff(OptimizationBarrier_31_io_y_eff),
    .io_y_c(OptimizationBarrier_31_io_y_c),
    .io_covSum(OptimizationBarrier_31_io_covSum),
    .metaAssert(OptimizationBarrier_31_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_32 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_32_io_x_ppn),
    .io_x_u(OptimizationBarrier_32_io_x_u),
    .io_x_ae(OptimizationBarrier_32_io_x_ae),
    .io_x_sw(OptimizationBarrier_32_io_x_sw),
    .io_x_sx(OptimizationBarrier_32_io_x_sx),
    .io_x_sr(OptimizationBarrier_32_io_x_sr),
    .io_x_pw(OptimizationBarrier_32_io_x_pw),
    .io_x_px(OptimizationBarrier_32_io_x_px),
    .io_x_pr(OptimizationBarrier_32_io_x_pr),
    .io_x_ppp(OptimizationBarrier_32_io_x_ppp),
    .io_x_pal(OptimizationBarrier_32_io_x_pal),
    .io_x_paa(OptimizationBarrier_32_io_x_paa),
    .io_x_eff(OptimizationBarrier_32_io_x_eff),
    .io_x_c(OptimizationBarrier_32_io_x_c),
    .io_y_ppn(OptimizationBarrier_32_io_y_ppn),
    .io_y_u(OptimizationBarrier_32_io_y_u),
    .io_y_ae(OptimizationBarrier_32_io_y_ae),
    .io_y_sw(OptimizationBarrier_32_io_y_sw),
    .io_y_sx(OptimizationBarrier_32_io_y_sx),
    .io_y_sr(OptimizationBarrier_32_io_y_sr),
    .io_y_pw(OptimizationBarrier_32_io_y_pw),
    .io_y_px(OptimizationBarrier_32_io_y_px),
    .io_y_pr(OptimizationBarrier_32_io_y_pr),
    .io_y_ppp(OptimizationBarrier_32_io_y_ppp),
    .io_y_pal(OptimizationBarrier_32_io_y_pal),
    .io_y_paa(OptimizationBarrier_32_io_y_paa),
    .io_y_eff(OptimizationBarrier_32_io_y_eff),
    .io_y_c(OptimizationBarrier_32_io_y_c),
    .io_covSum(OptimizationBarrier_32_io_covSum),
    .metaAssert(OptimizationBarrier_32_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_33 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_33_io_x_ppn),
    .io_x_u(OptimizationBarrier_33_io_x_u),
    .io_x_ae(OptimizationBarrier_33_io_x_ae),
    .io_x_sw(OptimizationBarrier_33_io_x_sw),
    .io_x_sx(OptimizationBarrier_33_io_x_sx),
    .io_x_sr(OptimizationBarrier_33_io_x_sr),
    .io_x_pw(OptimizationBarrier_33_io_x_pw),
    .io_x_px(OptimizationBarrier_33_io_x_px),
    .io_x_pr(OptimizationBarrier_33_io_x_pr),
    .io_x_ppp(OptimizationBarrier_33_io_x_ppp),
    .io_x_pal(OptimizationBarrier_33_io_x_pal),
    .io_x_paa(OptimizationBarrier_33_io_x_paa),
    .io_x_eff(OptimizationBarrier_33_io_x_eff),
    .io_x_c(OptimizationBarrier_33_io_x_c),
    .io_y_ppn(OptimizationBarrier_33_io_y_ppn),
    .io_y_u(OptimizationBarrier_33_io_y_u),
    .io_y_ae(OptimizationBarrier_33_io_y_ae),
    .io_y_sw(OptimizationBarrier_33_io_y_sw),
    .io_y_sx(OptimizationBarrier_33_io_y_sx),
    .io_y_sr(OptimizationBarrier_33_io_y_sr),
    .io_y_pw(OptimizationBarrier_33_io_y_pw),
    .io_y_px(OptimizationBarrier_33_io_y_px),
    .io_y_pr(OptimizationBarrier_33_io_y_pr),
    .io_y_ppp(OptimizationBarrier_33_io_y_ppp),
    .io_y_pal(OptimizationBarrier_33_io_y_pal),
    .io_y_paa(OptimizationBarrier_33_io_y_paa),
    .io_y_eff(OptimizationBarrier_33_io_y_eff),
    .io_y_c(OptimizationBarrier_33_io_y_c),
    .io_covSum(OptimizationBarrier_33_io_covSum),
    .metaAssert(OptimizationBarrier_33_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_34 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_34_io_x_ppn),
    .io_x_u(OptimizationBarrier_34_io_x_u),
    .io_x_ae(OptimizationBarrier_34_io_x_ae),
    .io_x_sw(OptimizationBarrier_34_io_x_sw),
    .io_x_sx(OptimizationBarrier_34_io_x_sx),
    .io_x_sr(OptimizationBarrier_34_io_x_sr),
    .io_x_pw(OptimizationBarrier_34_io_x_pw),
    .io_x_px(OptimizationBarrier_34_io_x_px),
    .io_x_pr(OptimizationBarrier_34_io_x_pr),
    .io_x_ppp(OptimizationBarrier_34_io_x_ppp),
    .io_x_pal(OptimizationBarrier_34_io_x_pal),
    .io_x_paa(OptimizationBarrier_34_io_x_paa),
    .io_x_eff(OptimizationBarrier_34_io_x_eff),
    .io_x_c(OptimizationBarrier_34_io_x_c),
    .io_y_ppn(OptimizationBarrier_34_io_y_ppn),
    .io_y_u(OptimizationBarrier_34_io_y_u),
    .io_y_ae(OptimizationBarrier_34_io_y_ae),
    .io_y_sw(OptimizationBarrier_34_io_y_sw),
    .io_y_sx(OptimizationBarrier_34_io_y_sx),
    .io_y_sr(OptimizationBarrier_34_io_y_sr),
    .io_y_pw(OptimizationBarrier_34_io_y_pw),
    .io_y_px(OptimizationBarrier_34_io_y_px),
    .io_y_pr(OptimizationBarrier_34_io_y_pr),
    .io_y_ppp(OptimizationBarrier_34_io_y_ppp),
    .io_y_pal(OptimizationBarrier_34_io_y_pal),
    .io_y_paa(OptimizationBarrier_34_io_y_paa),
    .io_y_eff(OptimizationBarrier_34_io_y_eff),
    .io_y_c(OptimizationBarrier_34_io_y_c),
    .io_covSum(OptimizationBarrier_34_io_covSum),
    .metaAssert(OptimizationBarrier_34_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_35 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_35_io_x_ppn),
    .io_x_u(OptimizationBarrier_35_io_x_u),
    .io_x_ae(OptimizationBarrier_35_io_x_ae),
    .io_x_sw(OptimizationBarrier_35_io_x_sw),
    .io_x_sx(OptimizationBarrier_35_io_x_sx),
    .io_x_sr(OptimizationBarrier_35_io_x_sr),
    .io_x_pw(OptimizationBarrier_35_io_x_pw),
    .io_x_px(OptimizationBarrier_35_io_x_px),
    .io_x_pr(OptimizationBarrier_35_io_x_pr),
    .io_x_ppp(OptimizationBarrier_35_io_x_ppp),
    .io_x_pal(OptimizationBarrier_35_io_x_pal),
    .io_x_paa(OptimizationBarrier_35_io_x_paa),
    .io_x_eff(OptimizationBarrier_35_io_x_eff),
    .io_x_c(OptimizationBarrier_35_io_x_c),
    .io_y_ppn(OptimizationBarrier_35_io_y_ppn),
    .io_y_u(OptimizationBarrier_35_io_y_u),
    .io_y_ae(OptimizationBarrier_35_io_y_ae),
    .io_y_sw(OptimizationBarrier_35_io_y_sw),
    .io_y_sx(OptimizationBarrier_35_io_y_sx),
    .io_y_sr(OptimizationBarrier_35_io_y_sr),
    .io_y_pw(OptimizationBarrier_35_io_y_pw),
    .io_y_px(OptimizationBarrier_35_io_y_px),
    .io_y_pr(OptimizationBarrier_35_io_y_pr),
    .io_y_ppp(OptimizationBarrier_35_io_y_ppp),
    .io_y_pal(OptimizationBarrier_35_io_y_pal),
    .io_y_paa(OptimizationBarrier_35_io_y_paa),
    .io_y_eff(OptimizationBarrier_35_io_y_eff),
    .io_y_c(OptimizationBarrier_35_io_y_c),
    .io_covSum(OptimizationBarrier_35_io_covSum),
    .metaAssert(OptimizationBarrier_35_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_36 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_36_io_x_ppn),
    .io_x_u(OptimizationBarrier_36_io_x_u),
    .io_x_ae(OptimizationBarrier_36_io_x_ae),
    .io_x_sw(OptimizationBarrier_36_io_x_sw),
    .io_x_sx(OptimizationBarrier_36_io_x_sx),
    .io_x_sr(OptimizationBarrier_36_io_x_sr),
    .io_x_pw(OptimizationBarrier_36_io_x_pw),
    .io_x_px(OptimizationBarrier_36_io_x_px),
    .io_x_pr(OptimizationBarrier_36_io_x_pr),
    .io_x_ppp(OptimizationBarrier_36_io_x_ppp),
    .io_x_pal(OptimizationBarrier_36_io_x_pal),
    .io_x_paa(OptimizationBarrier_36_io_x_paa),
    .io_x_eff(OptimizationBarrier_36_io_x_eff),
    .io_x_c(OptimizationBarrier_36_io_x_c),
    .io_y_ppn(OptimizationBarrier_36_io_y_ppn),
    .io_y_u(OptimizationBarrier_36_io_y_u),
    .io_y_ae(OptimizationBarrier_36_io_y_ae),
    .io_y_sw(OptimizationBarrier_36_io_y_sw),
    .io_y_sx(OptimizationBarrier_36_io_y_sx),
    .io_y_sr(OptimizationBarrier_36_io_y_sr),
    .io_y_pw(OptimizationBarrier_36_io_y_pw),
    .io_y_px(OptimizationBarrier_36_io_y_px),
    .io_y_pr(OptimizationBarrier_36_io_y_pr),
    .io_y_ppp(OptimizationBarrier_36_io_y_ppp),
    .io_y_pal(OptimizationBarrier_36_io_y_pal),
    .io_y_paa(OptimizationBarrier_36_io_y_paa),
    .io_y_eff(OptimizationBarrier_36_io_y_eff),
    .io_y_c(OptimizationBarrier_36_io_y_c),
    .io_covSum(OptimizationBarrier_36_io_covSum),
    .metaAssert(OptimizationBarrier_36_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_37 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_37_io_x_ppn),
    .io_x_u(OptimizationBarrier_37_io_x_u),
    .io_x_ae(OptimizationBarrier_37_io_x_ae),
    .io_x_sw(OptimizationBarrier_37_io_x_sw),
    .io_x_sx(OptimizationBarrier_37_io_x_sx),
    .io_x_sr(OptimizationBarrier_37_io_x_sr),
    .io_x_pw(OptimizationBarrier_37_io_x_pw),
    .io_x_px(OptimizationBarrier_37_io_x_px),
    .io_x_pr(OptimizationBarrier_37_io_x_pr),
    .io_x_ppp(OptimizationBarrier_37_io_x_ppp),
    .io_x_pal(OptimizationBarrier_37_io_x_pal),
    .io_x_paa(OptimizationBarrier_37_io_x_paa),
    .io_x_eff(OptimizationBarrier_37_io_x_eff),
    .io_x_c(OptimizationBarrier_37_io_x_c),
    .io_y_ppn(OptimizationBarrier_37_io_y_ppn),
    .io_y_u(OptimizationBarrier_37_io_y_u),
    .io_y_ae(OptimizationBarrier_37_io_y_ae),
    .io_y_sw(OptimizationBarrier_37_io_y_sw),
    .io_y_sx(OptimizationBarrier_37_io_y_sx),
    .io_y_sr(OptimizationBarrier_37_io_y_sr),
    .io_y_pw(OptimizationBarrier_37_io_y_pw),
    .io_y_px(OptimizationBarrier_37_io_y_px),
    .io_y_pr(OptimizationBarrier_37_io_y_pr),
    .io_y_ppp(OptimizationBarrier_37_io_y_ppp),
    .io_y_pal(OptimizationBarrier_37_io_y_pal),
    .io_y_paa(OptimizationBarrier_37_io_y_paa),
    .io_y_eff(OptimizationBarrier_37_io_y_eff),
    .io_y_c(OptimizationBarrier_37_io_y_c),
    .io_covSum(OptimizationBarrier_37_io_covSum),
    .metaAssert(OptimizationBarrier_37_metaAssert)
  );
  OptimizationBarrier OptimizationBarrier_38 ( // @[package.scala 236:25]
    .io_x_ppn(OptimizationBarrier_38_io_x_ppn),
    .io_x_u(OptimizationBarrier_38_io_x_u),
    .io_x_ae(OptimizationBarrier_38_io_x_ae),
    .io_x_sw(OptimizationBarrier_38_io_x_sw),
    .io_x_sx(OptimizationBarrier_38_io_x_sx),
    .io_x_sr(OptimizationBarrier_38_io_x_sr),
    .io_x_pw(OptimizationBarrier_38_io_x_pw),
    .io_x_px(OptimizationBarrier_38_io_x_px),
    .io_x_pr(OptimizationBarrier_38_io_x_pr),
    .io_x_ppp(OptimizationBarrier_38_io_x_ppp),
    .io_x_pal(OptimizationBarrier_38_io_x_pal),
    .io_x_paa(OptimizationBarrier_38_io_x_paa),
    .io_x_eff(OptimizationBarrier_38_io_x_eff),
    .io_x_c(OptimizationBarrier_38_io_x_c),
    .io_y_ppn(OptimizationBarrier_38_io_y_ppn),
    .io_y_u(OptimizationBarrier_38_io_y_u),
    .io_y_ae(OptimizationBarrier_38_io_y_ae),
    .io_y_sw(OptimizationBarrier_38_io_y_sw),
    .io_y_sx(OptimizationBarrier_38_io_y_sx),
    .io_y_sr(OptimizationBarrier_38_io_y_sr),
    .io_y_pw(OptimizationBarrier_38_io_y_pw),
    .io_y_px(OptimizationBarrier_38_io_y_px),
    .io_y_pr(OptimizationBarrier_38_io_y_pr),
    .io_y_ppp(OptimizationBarrier_38_io_y_ppp),
    .io_y_pal(OptimizationBarrier_38_io_y_pal),
    .io_y_paa(OptimizationBarrier_38_io_y_paa),
    .io_y_eff(OptimizationBarrier_38_io_y_eff),
    .io_y_c(OptimizationBarrier_38_io_y_c),
    .io_covSum(OptimizationBarrier_38_io_covSum),
    .metaAssert(OptimizationBarrier_38_metaAssert)
  );
  assign priv_s = io_ptw_status_prv[0]; // @[TLB.scala 177:20]
  assign priv_uses_vm = io_ptw_status_prv <= 2'h1; // @[TLB.scala 178:27]
  assign vm_enabled = io_ptw_ptbr_mode[3] & priv_uses_vm; // @[TLB.scala 179:83]
  assign vpn = io_req_bits_vaddr[38:12]; // @[TLB.scala 182:30]
  assign refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 183:44]
  assign _T_4 = state == 2'h1; // @[package.scala 15:47]
  assign _T_5 = state == 2'h3; // @[package.scala 15:47]
  assign _T_6 = _T_4 | _T_5; // @[package.scala 64:59]
  assign invalidate_refill = _T_6 | io_sfence_valid; // @[TLB.scala 185:88]
  assign _T_27 = special_entry_level < 2'h1; // @[TLB.scala 108:28]
  assign _T_29 = _T_27 ? vpn : 27'h0; // @[TLB.scala 109:28]
  assign _GEN_983 = {{7'd0}, OptimizationBarrier_io_y_ppn}; // @[TLB.scala 109:47]
  assign _T_30 = _T_29 | _GEN_983; // @[TLB.scala 109:47]
  assign _T_33 = special_entry_level < 2'h2; // @[TLB.scala 108:28]
  assign _T_35 = _T_33 ? vpn : 27'h0; // @[TLB.scala 109:28]
  assign _T_36 = _T_35 | _GEN_983; // @[TLB.scala 109:47]
  assign _T_38 = {OptimizationBarrier_io_y_ppn[19:18],_T_30[17:9],_T_36[8:0]}; // @[Cat.scala 29:58]
  assign _T_40 = vm_enabled ? {{8'd0}, _T_38} : io_req_bits_vaddr[39:12]; // @[TLB.scala 187:20]
  assign mpu_ppn = io_ptw_resp_valid ? {{8'd0}, refill_ppn} : _T_40; // @[TLB.scala 186:20]
  assign mpu_physaddr = {mpu_ppn,io_req_bits_vaddr[11:0]}; // @[Cat.scala 29:58]
  assign _T_44 = {io_ptw_status_debug,io_ptw_status_prv}; // @[Cat.scala 29:58]
  assign mpu_priv = io_ptw_resp_valid ? 3'h1 : _T_44; // @[TLB.scala 189:27]
  assign _T_45 = mpu_physaddr ^ 40'h3000; // @[Parameters.scala 137:31]
  assign _T_46 = {1'b0,$signed(_T_45)}; // @[Parameters.scala 137:49]
  assign _T_48 = $signed(_T_46) & -41'sh1000; // @[Parameters.scala 137:52]
  assign _T_49 = $signed(_T_48) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_50 = mpu_physaddr ^ 40'hc000000; // @[Parameters.scala 137:31]
  assign _T_51 = {1'b0,$signed(_T_50)}; // @[Parameters.scala 137:49]
  assign _T_53 = $signed(_T_51) & -41'sh4000000; // @[Parameters.scala 137:52]
  assign _T_54 = $signed(_T_53) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_55 = mpu_physaddr ^ 40'h2000000; // @[Parameters.scala 137:31]
  assign _T_56 = {1'b0,$signed(_T_55)}; // @[Parameters.scala 137:49]
  assign _T_58 = $signed(_T_56) & -41'sh10000; // @[Parameters.scala 137:52]
  assign _T_59 = $signed(_T_58) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_61 = {1'b0,$signed(mpu_physaddr)}; // @[Parameters.scala 137:49]
  assign _T_63 = $signed(_T_61) & -41'sh1000; // @[Parameters.scala 137:52]
  assign _T_64 = $signed(_T_63) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_65 = mpu_physaddr ^ 40'h10000; // @[Parameters.scala 137:31]
  assign _T_66 = {1'b0,$signed(_T_65)}; // @[Parameters.scala 137:49]
  assign _T_68 = $signed(_T_66) & -41'sh10000; // @[Parameters.scala 137:52]
  assign _T_69 = $signed(_T_68) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_70 = mpu_physaddr ^ 40'h80000000; // @[Parameters.scala 137:31]
  assign _T_71 = {1'b0,$signed(_T_70)}; // @[Parameters.scala 137:49]
  assign _T_73 = $signed(_T_71) & -41'sh10000000; // @[Parameters.scala 137:52]
  assign _T_74 = $signed(_T_73) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_75 = mpu_physaddr ^ 40'h60000000; // @[Parameters.scala 137:31]
  assign _T_76 = {1'b0,$signed(_T_75)}; // @[Parameters.scala 137:49]
  assign _T_78 = $signed(_T_76) & -41'sh20000000; // @[Parameters.scala 137:52]
  assign _T_79 = $signed(_T_78) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_81 = _T_49 | _T_54; // @[TLB.scala 195:67]
  assign _T_82 = _T_81 | _T_59; // @[TLB.scala 195:67]
  assign _T_83 = _T_82 | _T_64; // @[TLB.scala 195:67]
  assign _T_84 = _T_83 | _T_69; // @[TLB.scala 195:67]
  assign _T_85 = _T_84 | _T_74; // @[TLB.scala 195:67]
  assign legal_address = _T_85 | _T_79; // @[TLB.scala 195:67]
  assign _T_94 = $signed(_T_71) & 41'sh80000000; // @[Parameters.scala 137:52]
  assign _T_95 = $signed(_T_94) == 41'sh0; // @[Parameters.scala 137:67]
  assign cacheable = legal_address & _T_95; // @[TLB.scala 197:19]
  assign _T_155 = mpu_physaddr ^ 40'h8000000; // @[Parameters.scala 137:31]
  assign _T_156 = {1'b0,$signed(_T_155)}; // @[Parameters.scala 137:49]
  assign _T_158 = $signed(_T_156) & 41'shc8000000; // @[Parameters.scala 137:52]
  assign _T_159 = $signed(_T_158) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_172 = $signed(_T_61) & 41'shc8010000; // @[Parameters.scala 137:52]
  assign _T_173 = $signed(_T_172) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_180 = _T_173 | _T_159; // @[TLBPermissions.scala 82:66]
  assign _T_193 = mpu_priv <= 3'h3; // @[TLB.scala 200:39]
  assign deny_access_to_debug = _T_193 & _T_64; // @[TLB.scala 200:48]
  assign _T_206 = legal_address & ~deny_access_to_debug; // @[TLB.scala 201:41]
  assign prot_r = _T_206 & pmp_io_r; // @[TLB.scala 201:66]
  assign _T_217 = mpu_physaddr ^ 40'h40000000; // @[Parameters.scala 137:31]
  assign _T_218 = {1'b0,$signed(_T_217)}; // @[Parameters.scala 137:49]
  assign _T_220 = $signed(_T_218) & 41'shc0000000; // @[Parameters.scala 137:52]
  assign _T_221 = $signed(_T_220) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_225 = $signed(_T_71) & 41'shc0000000; // @[Parameters.scala 137:52]
  assign _T_226 = $signed(_T_225) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_228 = _T_180 | _T_221; // @[Parameters.scala 549:89]
  assign _T_229 = _T_228 | _T_226; // @[Parameters.scala 549:89]
  assign _T_239 = legal_address & _T_229; // @[TLB.scala 197:19]
  assign _T_241 = _T_239 & ~deny_access_to_debug; // @[TLB.scala 202:45]
  assign prot_w = _T_241 & pmp_io_w; // @[TLB.scala 202:70]
  assign prot_al = legal_address & _T_180; // @[TLB.scala 197:19]
  assign _T_341 = $signed(_T_61) & 41'shca000000; // @[Parameters.scala 137:52]
  assign _T_342 = $signed(_T_341) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_353 = _T_342 | _T_221; // @[Parameters.scala 549:89]
  assign _T_354 = _T_353 | _T_226; // @[Parameters.scala 549:89]
  assign _T_370 = legal_address & _T_354; // @[TLB.scala 197:19]
  assign _T_372 = _T_370 & ~deny_access_to_debug; // @[TLB.scala 206:40]
  assign prot_x = _T_372 & pmp_io_x; // @[TLB.scala 206:65]
  assign _T_393 = $signed(_T_61) & 41'shca012000; // @[Parameters.scala 137:52]
  assign _T_394 = $signed(_T_393) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_398 = $signed(_T_56) & 41'shca010000; // @[Parameters.scala 137:52]
  assign _T_399 = $signed(_T_398) == 41'sh0; // @[Parameters.scala 137:67]
  assign _T_410 = _T_394 | _T_399; // @[Parameters.scala 549:89]
  assign _T_411 = _T_410 | _T_159; // @[Parameters.scala 549:89]
  assign _T_412 = _T_411 | _T_221; // @[Parameters.scala 549:89]
  assign prot_eff = legal_address & _T_412; // @[TLB.scala 197:19]
  assign _T_417 = sectored_entries_0_valid_0 | sectored_entries_0_valid_1; // @[package.scala 64:59]
  assign _T_418 = _T_417 | sectored_entries_0_valid_2; // @[package.scala 64:59]
  assign _T_419 = _T_418 | sectored_entries_0_valid_3; // @[package.scala 64:59]
  assign _T_420 = sectored_entries_0_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_422 = _T_420[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_0 = _T_419 & _T_422; // @[TLB.scala 87:40]
  assign _T_423 = sectored_entries_1_valid_0 | sectored_entries_1_valid_1; // @[package.scala 64:59]
  assign _T_424 = _T_423 | sectored_entries_1_valid_2; // @[package.scala 64:59]
  assign _T_425 = _T_424 | sectored_entries_1_valid_3; // @[package.scala 64:59]
  assign _T_426 = sectored_entries_1_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_428 = _T_426[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_1 = _T_425 & _T_428; // @[TLB.scala 87:40]
  assign _T_429 = sectored_entries_2_valid_0 | sectored_entries_2_valid_1; // @[package.scala 64:59]
  assign _T_430 = _T_429 | sectored_entries_2_valid_2; // @[package.scala 64:59]
  assign _T_431 = _T_430 | sectored_entries_2_valid_3; // @[package.scala 64:59]
  assign _T_432 = sectored_entries_2_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_434 = _T_432[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_2 = _T_431 & _T_434; // @[TLB.scala 87:40]
  assign _T_435 = sectored_entries_3_valid_0 | sectored_entries_3_valid_1; // @[package.scala 64:59]
  assign _T_436 = _T_435 | sectored_entries_3_valid_2; // @[package.scala 64:59]
  assign _T_437 = _T_436 | sectored_entries_3_valid_3; // @[package.scala 64:59]
  assign _T_438 = sectored_entries_3_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_440 = _T_438[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_3 = _T_437 & _T_440; // @[TLB.scala 87:40]
  assign _T_441 = sectored_entries_4_valid_0 | sectored_entries_4_valid_1; // @[package.scala 64:59]
  assign _T_442 = _T_441 | sectored_entries_4_valid_2; // @[package.scala 64:59]
  assign _T_443 = _T_442 | sectored_entries_4_valid_3; // @[package.scala 64:59]
  assign _T_444 = sectored_entries_4_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_446 = _T_444[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_4 = _T_443 & _T_446; // @[TLB.scala 87:40]
  assign _T_447 = sectored_entries_5_valid_0 | sectored_entries_5_valid_1; // @[package.scala 64:59]
  assign _T_448 = _T_447 | sectored_entries_5_valid_2; // @[package.scala 64:59]
  assign _T_449 = _T_448 | sectored_entries_5_valid_3; // @[package.scala 64:59]
  assign _T_450 = sectored_entries_5_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_452 = _T_450[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_5 = _T_449 & _T_452; // @[TLB.scala 87:40]
  assign _T_453 = sectored_entries_6_valid_0 | sectored_entries_6_valid_1; // @[package.scala 64:59]
  assign _T_454 = _T_453 | sectored_entries_6_valid_2; // @[package.scala 64:59]
  assign _T_455 = _T_454 | sectored_entries_6_valid_3; // @[package.scala 64:59]
  assign _T_456 = sectored_entries_6_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_458 = _T_456[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_6 = _T_455 & _T_458; // @[TLB.scala 87:40]
  assign _T_459 = sectored_entries_7_valid_0 | sectored_entries_7_valid_1; // @[package.scala 64:59]
  assign _T_460 = _T_459 | sectored_entries_7_valid_2; // @[package.scala 64:59]
  assign _T_461 = _T_460 | sectored_entries_7_valid_3; // @[package.scala 64:59]
  assign _T_462 = sectored_entries_7_tag ^ vpn; // @[TLB.scala 88:41]
  assign _T_464 = _T_462[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_7 = _T_461 & _T_464; // @[TLB.scala 87:40]
  assign _T_469 = superpage_entries_0_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _T_471 = superpage_entries_0_valid_0 & _T_469; // @[TLB.scala 95:29]
  assign _T_472 = superpage_entries_0_level < 2'h1; // @[TLB.scala 94:28]
  assign _T_476 = superpage_entries_0_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _T_477 = _T_472 | _T_476; // @[TLB.scala 95:40]
  assign superpage_hits_0 = _T_471 & _T_477; // @[TLB.scala 95:29]
  assign _T_489 = superpage_entries_1_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _T_491 = superpage_entries_1_valid_0 & _T_489; // @[TLB.scala 95:29]
  assign _T_492 = superpage_entries_1_level < 2'h1; // @[TLB.scala 94:28]
  assign _T_496 = superpage_entries_1_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _T_497 = _T_492 | _T_496; // @[TLB.scala 95:40]
  assign superpage_hits_1 = _T_491 & _T_497; // @[TLB.scala 95:29]
  assign _T_509 = superpage_entries_2_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _T_511 = superpage_entries_2_valid_0 & _T_509; // @[TLB.scala 95:29]
  assign _T_512 = superpage_entries_2_level < 2'h1; // @[TLB.scala 94:28]
  assign _T_516 = superpage_entries_2_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _T_517 = _T_512 | _T_516; // @[TLB.scala 95:40]
  assign superpage_hits_2 = _T_511 & _T_517; // @[TLB.scala 95:29]
  assign _T_529 = superpage_entries_3_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _T_531 = superpage_entries_3_valid_0 & _T_529; // @[TLB.scala 95:29]
  assign _T_532 = superpage_entries_3_level < 2'h1; // @[TLB.scala 94:28]
  assign _T_536 = superpage_entries_3_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _T_537 = _T_532 | _T_536; // @[TLB.scala 95:40]
  assign superpage_hits_3 = _T_531 & _T_537; // @[TLB.scala 95:29]
  assign _GEN_1 = 2'h1 == vpn[1:0] ? sectored_entries_0_valid_1 : sectored_entries_0_valid_0; // @[TLB.scala 100:18]
  assign _GEN_2 = 2'h2 == vpn[1:0] ? sectored_entries_0_valid_2 : _GEN_1; // @[TLB.scala 100:18]
  assign _GEN_3 = 2'h3 == vpn[1:0] ? sectored_entries_0_valid_3 : _GEN_2; // @[TLB.scala 100:18]
  assign _T_549 = _GEN_3 & _T_422; // @[TLB.scala 100:18]
  assign hitsVec_0 = vm_enabled & _T_549; // @[TLB.scala 211:44]
  assign _GEN_5 = 2'h1 == vpn[1:0] ? sectored_entries_1_valid_1 : sectored_entries_1_valid_0; // @[TLB.scala 100:18]
  assign _GEN_6 = 2'h2 == vpn[1:0] ? sectored_entries_1_valid_2 : _GEN_5; // @[TLB.scala 100:18]
  assign _GEN_7 = 2'h3 == vpn[1:0] ? sectored_entries_1_valid_3 : _GEN_6; // @[TLB.scala 100:18]
  assign _T_554 = _GEN_7 & _T_428; // @[TLB.scala 100:18]
  assign hitsVec_1 = vm_enabled & _T_554; // @[TLB.scala 211:44]
  assign _GEN_9 = 2'h1 == vpn[1:0] ? sectored_entries_2_valid_1 : sectored_entries_2_valid_0; // @[TLB.scala 100:18]
  assign _GEN_10 = 2'h2 == vpn[1:0] ? sectored_entries_2_valid_2 : _GEN_9; // @[TLB.scala 100:18]
  assign _GEN_11 = 2'h3 == vpn[1:0] ? sectored_entries_2_valid_3 : _GEN_10; // @[TLB.scala 100:18]
  assign _T_559 = _GEN_11 & _T_434; // @[TLB.scala 100:18]
  assign hitsVec_2 = vm_enabled & _T_559; // @[TLB.scala 211:44]
  assign _GEN_13 = 2'h1 == vpn[1:0] ? sectored_entries_3_valid_1 : sectored_entries_3_valid_0; // @[TLB.scala 100:18]
  assign _GEN_14 = 2'h2 == vpn[1:0] ? sectored_entries_3_valid_2 : _GEN_13; // @[TLB.scala 100:18]
  assign _GEN_15 = 2'h3 == vpn[1:0] ? sectored_entries_3_valid_3 : _GEN_14; // @[TLB.scala 100:18]
  assign _T_564 = _GEN_15 & _T_440; // @[TLB.scala 100:18]
  assign hitsVec_3 = vm_enabled & _T_564; // @[TLB.scala 211:44]
  assign _GEN_17 = 2'h1 == vpn[1:0] ? sectored_entries_4_valid_1 : sectored_entries_4_valid_0; // @[TLB.scala 100:18]
  assign _GEN_18 = 2'h2 == vpn[1:0] ? sectored_entries_4_valid_2 : _GEN_17; // @[TLB.scala 100:18]
  assign _GEN_19 = 2'h3 == vpn[1:0] ? sectored_entries_4_valid_3 : _GEN_18; // @[TLB.scala 100:18]
  assign _T_569 = _GEN_19 & _T_446; // @[TLB.scala 100:18]
  assign hitsVec_4 = vm_enabled & _T_569; // @[TLB.scala 211:44]
  assign _GEN_21 = 2'h1 == vpn[1:0] ? sectored_entries_5_valid_1 : sectored_entries_5_valid_0; // @[TLB.scala 100:18]
  assign _GEN_22 = 2'h2 == vpn[1:0] ? sectored_entries_5_valid_2 : _GEN_21; // @[TLB.scala 100:18]
  assign _GEN_23 = 2'h3 == vpn[1:0] ? sectored_entries_5_valid_3 : _GEN_22; // @[TLB.scala 100:18]
  assign _T_574 = _GEN_23 & _T_452; // @[TLB.scala 100:18]
  assign hitsVec_5 = vm_enabled & _T_574; // @[TLB.scala 211:44]
  assign _GEN_25 = 2'h1 == vpn[1:0] ? sectored_entries_6_valid_1 : sectored_entries_6_valid_0; // @[TLB.scala 100:18]
  assign _GEN_26 = 2'h2 == vpn[1:0] ? sectored_entries_6_valid_2 : _GEN_25; // @[TLB.scala 100:18]
  assign _GEN_27 = 2'h3 == vpn[1:0] ? sectored_entries_6_valid_3 : _GEN_26; // @[TLB.scala 100:18]
  assign _T_579 = _GEN_27 & _T_458; // @[TLB.scala 100:18]
  assign hitsVec_6 = vm_enabled & _T_579; // @[TLB.scala 211:44]
  assign _GEN_29 = 2'h1 == vpn[1:0] ? sectored_entries_7_valid_1 : sectored_entries_7_valid_0; // @[TLB.scala 100:18]
  assign _GEN_30 = 2'h2 == vpn[1:0] ? sectored_entries_7_valid_2 : _GEN_29; // @[TLB.scala 100:18]
  assign _GEN_31 = 2'h3 == vpn[1:0] ? sectored_entries_7_valid_3 : _GEN_30; // @[TLB.scala 100:18]
  assign _T_584 = _GEN_31 & _T_464; // @[TLB.scala 100:18]
  assign hitsVec_7 = vm_enabled & _T_584; // @[TLB.scala 211:44]
  assign hitsVec_8 = vm_enabled & superpage_hits_0; // @[TLB.scala 211:44]
  assign hitsVec_9 = vm_enabled & superpage_hits_1; // @[TLB.scala 211:44]
  assign hitsVec_10 = vm_enabled & superpage_hits_2; // @[TLB.scala 211:44]
  assign hitsVec_11 = vm_enabled & superpage_hits_3; // @[TLB.scala 211:44]
  assign _T_673 = special_entry_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _T_675 = special_entry_valid_0 & _T_673; // @[TLB.scala 95:29]
  assign _T_680 = special_entry_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _T_681 = _T_27 | _T_680; // @[TLB.scala 95:40]
  assign _T_682 = _T_675 & _T_681; // @[TLB.scala 95:29]
  assign _T_687 = special_entry_tag[8:0] == vpn[8:0]; // @[TLB.scala 95:77]
  assign _T_688 = _T_33 | _T_687; // @[TLB.scala 95:40]
  assign _T_689 = _T_682 & _T_688; // @[TLB.scala 95:29]
  assign hitsVec_12 = vm_enabled & _T_689; // @[TLB.scala 211:44]
  assign _T_694 = {hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[Cat.scala 29:58]
  assign real_hits = {hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_694}; // @[Cat.scala 29:58]
  assign hits = {~vm_enabled,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_694}; // @[Cat.scala 29:58]
  assign _GEN_33 = 2'h1 == vpn[1:0] ? sectored_entries_0_data_1 : sectored_entries_0_data_0;
  assign _GEN_34 = 2'h2 == vpn[1:0] ? sectored_entries_0_data_2 : _GEN_33;
  assign _GEN_35 = 2'h3 == vpn[1:0] ? sectored_entries_0_data_3 : _GEN_34;
  assign _GEN_37 = 2'h1 == vpn[1:0] ? sectored_entries_1_data_1 : sectored_entries_1_data_0;
  assign _GEN_38 = 2'h2 == vpn[1:0] ? sectored_entries_1_data_2 : _GEN_37;
  assign _GEN_39 = 2'h3 == vpn[1:0] ? sectored_entries_1_data_3 : _GEN_38;
  assign _GEN_41 = 2'h1 == vpn[1:0] ? sectored_entries_2_data_1 : sectored_entries_2_data_0;
  assign _GEN_42 = 2'h2 == vpn[1:0] ? sectored_entries_2_data_2 : _GEN_41;
  assign _GEN_43 = 2'h3 == vpn[1:0] ? sectored_entries_2_data_3 : _GEN_42;
  assign _GEN_45 = 2'h1 == vpn[1:0] ? sectored_entries_3_data_1 : sectored_entries_3_data_0;
  assign _GEN_46 = 2'h2 == vpn[1:0] ? sectored_entries_3_data_2 : _GEN_45;
  assign _GEN_47 = 2'h3 == vpn[1:0] ? sectored_entries_3_data_3 : _GEN_46;
  assign _GEN_49 = 2'h1 == vpn[1:0] ? sectored_entries_4_data_1 : sectored_entries_4_data_0;
  assign _GEN_50 = 2'h2 == vpn[1:0] ? sectored_entries_4_data_2 : _GEN_49;
  assign _GEN_51 = 2'h3 == vpn[1:0] ? sectored_entries_4_data_3 : _GEN_50;
  assign _GEN_53 = 2'h1 == vpn[1:0] ? sectored_entries_5_data_1 : sectored_entries_5_data_0;
  assign _GEN_54 = 2'h2 == vpn[1:0] ? sectored_entries_5_data_2 : _GEN_53;
  assign _GEN_55 = 2'h3 == vpn[1:0] ? sectored_entries_5_data_3 : _GEN_54;
  assign _GEN_57 = 2'h1 == vpn[1:0] ? sectored_entries_6_data_1 : sectored_entries_6_data_0;
  assign _GEN_58 = 2'h2 == vpn[1:0] ? sectored_entries_6_data_2 : _GEN_57;
  assign _GEN_59 = 2'h3 == vpn[1:0] ? sectored_entries_6_data_3 : _GEN_58;
  assign _GEN_61 = 2'h1 == vpn[1:0] ? sectored_entries_7_data_1 : sectored_entries_7_data_0;
  assign _GEN_62 = 2'h2 == vpn[1:0] ? sectored_entries_7_data_2 : _GEN_61;
  assign _GEN_63 = 2'h3 == vpn[1:0] ? sectored_entries_7_data_3 : _GEN_62;
  assign _T_876 = _T_472 ? vpn : 27'h0; // @[TLB.scala 109:28]
  assign _GEN_985 = {{7'd0}, OptimizationBarrier_9_io_y_ppn}; // @[TLB.scala 109:47]
  assign _T_877 = _T_876 | _GEN_985; // @[TLB.scala 109:47]
  assign _T_883 = vpn | _GEN_985; // @[TLB.scala 109:47]
  assign _T_885 = {OptimizationBarrier_9_io_y_ppn[19:18],_T_877[17:9],_T_883[8:0]}; // @[Cat.scala 29:58]
  assign _T_907 = _T_492 ? vpn : 27'h0; // @[TLB.scala 109:28]
  assign _GEN_987 = {{7'd0}, OptimizationBarrier_10_io_y_ppn}; // @[TLB.scala 109:47]
  assign _T_908 = _T_907 | _GEN_987; // @[TLB.scala 109:47]
  assign _T_914 = vpn | _GEN_987; // @[TLB.scala 109:47]
  assign _T_916 = {OptimizationBarrier_10_io_y_ppn[19:18],_T_908[17:9],_T_914[8:0]}; // @[Cat.scala 29:58]
  assign _T_938 = _T_512 ? vpn : 27'h0; // @[TLB.scala 109:28]
  assign _GEN_989 = {{7'd0}, OptimizationBarrier_11_io_y_ppn}; // @[TLB.scala 109:47]
  assign _T_939 = _T_938 | _GEN_989; // @[TLB.scala 109:47]
  assign _T_945 = vpn | _GEN_989; // @[TLB.scala 109:47]
  assign _T_947 = {OptimizationBarrier_11_io_y_ppn[19:18],_T_939[17:9],_T_945[8:0]}; // @[Cat.scala 29:58]
  assign _T_969 = _T_532 ? vpn : 27'h0; // @[TLB.scala 109:28]
  assign _GEN_991 = {{7'd0}, OptimizationBarrier_12_io_y_ppn}; // @[TLB.scala 109:47]
  assign _T_970 = _T_969 | _GEN_991; // @[TLB.scala 109:47]
  assign _T_976 = vpn | _GEN_991; // @[TLB.scala 109:47]
  assign _T_978 = {OptimizationBarrier_12_io_y_ppn[19:18],_T_970[17:9],_T_976[8:0]}; // @[Cat.scala 29:58]
  assign _GEN_993 = {{7'd0}, OptimizationBarrier_13_io_y_ppn}; // @[TLB.scala 109:47]
  assign _T_1001 = _T_29 | _GEN_993; // @[TLB.scala 109:47]
  assign _T_1007 = _T_35 | _GEN_993; // @[TLB.scala 109:47]
  assign _T_1009 = {OptimizationBarrier_13_io_y_ppn[19:18],_T_1001[17:9],_T_1007[8:0]}; // @[Cat.scala 29:58]
  assign _T_1011 = hitsVec_0 ? OptimizationBarrier_1_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1012 = hitsVec_1 ? OptimizationBarrier_2_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1013 = hitsVec_2 ? OptimizationBarrier_3_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1014 = hitsVec_3 ? OptimizationBarrier_4_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1015 = hitsVec_4 ? OptimizationBarrier_5_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1016 = hitsVec_5 ? OptimizationBarrier_6_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1017 = hitsVec_6 ? OptimizationBarrier_7_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1018 = hitsVec_7 ? OptimizationBarrier_8_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _T_1019 = hitsVec_8 ? _T_885 : 20'h0; // @[Mux.scala 27:72]
  assign _T_1020 = hitsVec_9 ? _T_916 : 20'h0; // @[Mux.scala 27:72]
  assign _T_1021 = hitsVec_10 ? _T_947 : 20'h0; // @[Mux.scala 27:72]
  assign _T_1022 = hitsVec_11 ? _T_978 : 20'h0; // @[Mux.scala 27:72]
  assign _T_1023 = hitsVec_12 ? _T_1009 : 20'h0; // @[Mux.scala 27:72]
  assign _T_1024 = vm_enabled ? 20'h0 : vpn[19:0]; // @[Mux.scala 27:72]
  assign _T_1025 = _T_1011 | _T_1012; // @[Mux.scala 27:72]
  assign _T_1026 = _T_1025 | _T_1013; // @[Mux.scala 27:72]
  assign _T_1027 = _T_1026 | _T_1014; // @[Mux.scala 27:72]
  assign _T_1028 = _T_1027 | _T_1015; // @[Mux.scala 27:72]
  assign _T_1029 = _T_1028 | _T_1016; // @[Mux.scala 27:72]
  assign _T_1030 = _T_1029 | _T_1017; // @[Mux.scala 27:72]
  assign _T_1031 = _T_1030 | _T_1018; // @[Mux.scala 27:72]
  assign _T_1032 = _T_1031 | _T_1019; // @[Mux.scala 27:72]
  assign _T_1033 = _T_1032 | _T_1020; // @[Mux.scala 27:72]
  assign _T_1034 = _T_1033 | _T_1021; // @[Mux.scala 27:72]
  assign _T_1035 = _T_1034 | _T_1022; // @[Mux.scala 27:72]
  assign _T_1036 = _T_1035 | _T_1023; // @[Mux.scala 27:72]
  assign ppn = _T_1036 | _T_1024; // @[Mux.scala 27:72]
  assign _T_1039 = io_ptw_resp_bits_pte_g & io_ptw_resp_bits_pte_v; // @[TLB.scala 223:25]
  assign _T_1041 = io_ptw_resp_bits_pte_x & ~io_ptw_resp_bits_pte_w; // @[PTW.scala 69:44]
  assign _T_1042 = io_ptw_resp_bits_pte_r | _T_1041; // @[PTW.scala 69:38]
  assign _T_1043 = io_ptw_resp_bits_pte_v & _T_1042; // @[PTW.scala 69:32]
  assign _T_1044 = _T_1043 & io_ptw_resp_bits_pte_a; // @[PTW.scala 69:52]
  assign _T_1045 = _T_1044 & io_ptw_resp_bits_pte_r; // @[PTW.scala 73:35]
  assign _T_1051 = _T_1044 & io_ptw_resp_bits_pte_w; // @[PTW.scala 74:35]
  assign _T_1052 = _T_1051 & io_ptw_resp_bits_pte_d; // @[PTW.scala 74:40]
  assign _T_1058 = _T_1044 & io_ptw_resp_bits_pte_x; // @[PTW.scala 75:35]
  assign _T_1068 = {prot_x,prot_r,_T_239,prot_al,prot_al,prot_eff,cacheable,1'h0}; // @[TLB.scala 123:24]
  assign _T_1076 = {refill_ppn,io_ptw_resp_bits_pte_u,_T_1039,io_ptw_resp_bits_ae,_T_1052,_T_1058,_T_1045,prot_w,_T_1068}; // @[TLB.scala 123:24]
  assign _GEN_64 = invalidate_refill ? 1'h0 : 1'h1; // @[TLB.scala 240:34]
  assign _T_1077 = io_ptw_resp_bits_level < 2'h2; // @[TLB.scala 242:40]
  assign _T_1078 = r_superpage_repl_addr == 2'h0; // @[TLB.scala 243:82]
  assign _GEN_67 = _T_1078 ? _GEN_64 : superpage_entries_0_valid_0; // @[TLB.scala 243:89]
  assign _T_1095 = r_superpage_repl_addr == 2'h1; // @[TLB.scala 243:82]
  assign _GEN_71 = _T_1095 ? _GEN_64 : superpage_entries_1_valid_0; // @[TLB.scala 243:89]
  assign _T_1112 = r_superpage_repl_addr == 2'h2; // @[TLB.scala 243:82]
  assign _GEN_75 = _T_1112 ? _GEN_64 : superpage_entries_2_valid_0; // @[TLB.scala 243:89]
  assign _T_1129 = r_superpage_repl_addr == 2'h3; // @[TLB.scala 243:82]
  assign _GEN_79 = _T_1129 ? _GEN_64 : superpage_entries_3_valid_0; // @[TLB.scala 243:89]
  assign _T_1146 = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; // @[TLB.scala 248:22]
  assign _T_1147 = _T_1146 == 3'h0; // @[TLB.scala 249:65]
  assign _GEN_81 = r_sectored_hit ? sectored_entries_0_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_82 = r_sectored_hit ? sectored_entries_0_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_83 = r_sectored_hit ? sectored_entries_0_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_84 = r_sectored_hit ? sectored_entries_0_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_995 = 2'h0 == r_refill_tag[1:0]; // @[TLB.scala 122:16]
  assign _GEN_85 = _GEN_995 | _GEN_81; // @[TLB.scala 122:16]
  assign _GEN_996 = 2'h1 == r_refill_tag[1:0]; // @[TLB.scala 122:16]
  assign _GEN_86 = _GEN_996 | _GEN_82; // @[TLB.scala 122:16]
  assign _GEN_997 = 2'h2 == r_refill_tag[1:0]; // @[TLB.scala 122:16]
  assign _GEN_87 = _GEN_997 | _GEN_83; // @[TLB.scala 122:16]
  assign _GEN_998 = 2'h3 == r_refill_tag[1:0]; // @[TLB.scala 122:16]
  assign _GEN_88 = _GEN_998 | _GEN_84; // @[TLB.scala 122:16]
  assign _GEN_93 = invalidate_refill ? 1'h0 : _GEN_85; // @[TLB.scala 252:34]
  assign _GEN_94 = invalidate_refill ? 1'h0 : _GEN_86; // @[TLB.scala 252:34]
  assign _GEN_95 = invalidate_refill ? 1'h0 : _GEN_87; // @[TLB.scala 252:34]
  assign _GEN_96 = invalidate_refill ? 1'h0 : _GEN_88; // @[TLB.scala 252:34]
  assign _GEN_97 = _T_1147 ? _GEN_93 : sectored_entries_0_valid_0; // @[TLB.scala 249:72]
  assign _GEN_98 = _T_1147 ? _GEN_94 : sectored_entries_0_valid_1; // @[TLB.scala 249:72]
  assign _GEN_99 = _T_1147 ? _GEN_95 : sectored_entries_0_valid_2; // @[TLB.scala 249:72]
  assign _GEN_100 = _T_1147 ? _GEN_96 : sectored_entries_0_valid_3; // @[TLB.scala 249:72]
  assign _T_1165 = _T_1146 == 3'h1; // @[TLB.scala 249:65]
  assign _GEN_107 = r_sectored_hit ? sectored_entries_1_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_108 = r_sectored_hit ? sectored_entries_1_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_109 = r_sectored_hit ? sectored_entries_1_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_110 = r_sectored_hit ? sectored_entries_1_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_111 = _GEN_995 | _GEN_107; // @[TLB.scala 122:16]
  assign _GEN_112 = _GEN_996 | _GEN_108; // @[TLB.scala 122:16]
  assign _GEN_113 = _GEN_997 | _GEN_109; // @[TLB.scala 122:16]
  assign _GEN_114 = _GEN_998 | _GEN_110; // @[TLB.scala 122:16]
  assign _GEN_119 = invalidate_refill ? 1'h0 : _GEN_111; // @[TLB.scala 252:34]
  assign _GEN_120 = invalidate_refill ? 1'h0 : _GEN_112; // @[TLB.scala 252:34]
  assign _GEN_121 = invalidate_refill ? 1'h0 : _GEN_113; // @[TLB.scala 252:34]
  assign _GEN_122 = invalidate_refill ? 1'h0 : _GEN_114; // @[TLB.scala 252:34]
  assign _GEN_123 = _T_1165 ? _GEN_119 : sectored_entries_1_valid_0; // @[TLB.scala 249:72]
  assign _GEN_124 = _T_1165 ? _GEN_120 : sectored_entries_1_valid_1; // @[TLB.scala 249:72]
  assign _GEN_125 = _T_1165 ? _GEN_121 : sectored_entries_1_valid_2; // @[TLB.scala 249:72]
  assign _GEN_126 = _T_1165 ? _GEN_122 : sectored_entries_1_valid_3; // @[TLB.scala 249:72]
  assign _T_1183 = _T_1146 == 3'h2; // @[TLB.scala 249:65]
  assign _GEN_133 = r_sectored_hit ? sectored_entries_2_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_134 = r_sectored_hit ? sectored_entries_2_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_135 = r_sectored_hit ? sectored_entries_2_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_136 = r_sectored_hit ? sectored_entries_2_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_137 = _GEN_995 | _GEN_133; // @[TLB.scala 122:16]
  assign _GEN_138 = _GEN_996 | _GEN_134; // @[TLB.scala 122:16]
  assign _GEN_139 = _GEN_997 | _GEN_135; // @[TLB.scala 122:16]
  assign _GEN_140 = _GEN_998 | _GEN_136; // @[TLB.scala 122:16]
  assign _GEN_145 = invalidate_refill ? 1'h0 : _GEN_137; // @[TLB.scala 252:34]
  assign _GEN_146 = invalidate_refill ? 1'h0 : _GEN_138; // @[TLB.scala 252:34]
  assign _GEN_147 = invalidate_refill ? 1'h0 : _GEN_139; // @[TLB.scala 252:34]
  assign _GEN_148 = invalidate_refill ? 1'h0 : _GEN_140; // @[TLB.scala 252:34]
  assign _GEN_149 = _T_1183 ? _GEN_145 : sectored_entries_2_valid_0; // @[TLB.scala 249:72]
  assign _GEN_150 = _T_1183 ? _GEN_146 : sectored_entries_2_valid_1; // @[TLB.scala 249:72]
  assign _GEN_151 = _T_1183 ? _GEN_147 : sectored_entries_2_valid_2; // @[TLB.scala 249:72]
  assign _GEN_152 = _T_1183 ? _GEN_148 : sectored_entries_2_valid_3; // @[TLB.scala 249:72]
  assign _T_1201 = _T_1146 == 3'h3; // @[TLB.scala 249:65]
  assign _GEN_159 = r_sectored_hit ? sectored_entries_3_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_160 = r_sectored_hit ? sectored_entries_3_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_161 = r_sectored_hit ? sectored_entries_3_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_162 = r_sectored_hit ? sectored_entries_3_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_163 = _GEN_995 | _GEN_159; // @[TLB.scala 122:16]
  assign _GEN_164 = _GEN_996 | _GEN_160; // @[TLB.scala 122:16]
  assign _GEN_165 = _GEN_997 | _GEN_161; // @[TLB.scala 122:16]
  assign _GEN_166 = _GEN_998 | _GEN_162; // @[TLB.scala 122:16]
  assign _GEN_171 = invalidate_refill ? 1'h0 : _GEN_163; // @[TLB.scala 252:34]
  assign _GEN_172 = invalidate_refill ? 1'h0 : _GEN_164; // @[TLB.scala 252:34]
  assign _GEN_173 = invalidate_refill ? 1'h0 : _GEN_165; // @[TLB.scala 252:34]
  assign _GEN_174 = invalidate_refill ? 1'h0 : _GEN_166; // @[TLB.scala 252:34]
  assign _GEN_175 = _T_1201 ? _GEN_171 : sectored_entries_3_valid_0; // @[TLB.scala 249:72]
  assign _GEN_176 = _T_1201 ? _GEN_172 : sectored_entries_3_valid_1; // @[TLB.scala 249:72]
  assign _GEN_177 = _T_1201 ? _GEN_173 : sectored_entries_3_valid_2; // @[TLB.scala 249:72]
  assign _GEN_178 = _T_1201 ? _GEN_174 : sectored_entries_3_valid_3; // @[TLB.scala 249:72]
  assign _T_1219 = _T_1146 == 3'h4; // @[TLB.scala 249:65]
  assign _GEN_185 = r_sectored_hit ? sectored_entries_4_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_186 = r_sectored_hit ? sectored_entries_4_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_187 = r_sectored_hit ? sectored_entries_4_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_188 = r_sectored_hit ? sectored_entries_4_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_189 = _GEN_995 | _GEN_185; // @[TLB.scala 122:16]
  assign _GEN_190 = _GEN_996 | _GEN_186; // @[TLB.scala 122:16]
  assign _GEN_191 = _GEN_997 | _GEN_187; // @[TLB.scala 122:16]
  assign _GEN_192 = _GEN_998 | _GEN_188; // @[TLB.scala 122:16]
  assign _GEN_197 = invalidate_refill ? 1'h0 : _GEN_189; // @[TLB.scala 252:34]
  assign _GEN_198 = invalidate_refill ? 1'h0 : _GEN_190; // @[TLB.scala 252:34]
  assign _GEN_199 = invalidate_refill ? 1'h0 : _GEN_191; // @[TLB.scala 252:34]
  assign _GEN_200 = invalidate_refill ? 1'h0 : _GEN_192; // @[TLB.scala 252:34]
  assign _GEN_201 = _T_1219 ? _GEN_197 : sectored_entries_4_valid_0; // @[TLB.scala 249:72]
  assign _GEN_202 = _T_1219 ? _GEN_198 : sectored_entries_4_valid_1; // @[TLB.scala 249:72]
  assign _GEN_203 = _T_1219 ? _GEN_199 : sectored_entries_4_valid_2; // @[TLB.scala 249:72]
  assign _GEN_204 = _T_1219 ? _GEN_200 : sectored_entries_4_valid_3; // @[TLB.scala 249:72]
  assign _T_1237 = _T_1146 == 3'h5; // @[TLB.scala 249:65]
  assign _GEN_211 = r_sectored_hit ? sectored_entries_5_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_212 = r_sectored_hit ? sectored_entries_5_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_213 = r_sectored_hit ? sectored_entries_5_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_214 = r_sectored_hit ? sectored_entries_5_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_215 = _GEN_995 | _GEN_211; // @[TLB.scala 122:16]
  assign _GEN_216 = _GEN_996 | _GEN_212; // @[TLB.scala 122:16]
  assign _GEN_217 = _GEN_997 | _GEN_213; // @[TLB.scala 122:16]
  assign _GEN_218 = _GEN_998 | _GEN_214; // @[TLB.scala 122:16]
  assign _GEN_223 = invalidate_refill ? 1'h0 : _GEN_215; // @[TLB.scala 252:34]
  assign _GEN_224 = invalidate_refill ? 1'h0 : _GEN_216; // @[TLB.scala 252:34]
  assign _GEN_225 = invalidate_refill ? 1'h0 : _GEN_217; // @[TLB.scala 252:34]
  assign _GEN_226 = invalidate_refill ? 1'h0 : _GEN_218; // @[TLB.scala 252:34]
  assign _GEN_227 = _T_1237 ? _GEN_223 : sectored_entries_5_valid_0; // @[TLB.scala 249:72]
  assign _GEN_228 = _T_1237 ? _GEN_224 : sectored_entries_5_valid_1; // @[TLB.scala 249:72]
  assign _GEN_229 = _T_1237 ? _GEN_225 : sectored_entries_5_valid_2; // @[TLB.scala 249:72]
  assign _GEN_230 = _T_1237 ? _GEN_226 : sectored_entries_5_valid_3; // @[TLB.scala 249:72]
  assign _T_1255 = _T_1146 == 3'h6; // @[TLB.scala 249:65]
  assign _GEN_237 = r_sectored_hit ? sectored_entries_6_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_238 = r_sectored_hit ? sectored_entries_6_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_239 = r_sectored_hit ? sectored_entries_6_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_240 = r_sectored_hit ? sectored_entries_6_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_241 = _GEN_995 | _GEN_237; // @[TLB.scala 122:16]
  assign _GEN_242 = _GEN_996 | _GEN_238; // @[TLB.scala 122:16]
  assign _GEN_243 = _GEN_997 | _GEN_239; // @[TLB.scala 122:16]
  assign _GEN_244 = _GEN_998 | _GEN_240; // @[TLB.scala 122:16]
  assign _GEN_249 = invalidate_refill ? 1'h0 : _GEN_241; // @[TLB.scala 252:34]
  assign _GEN_250 = invalidate_refill ? 1'h0 : _GEN_242; // @[TLB.scala 252:34]
  assign _GEN_251 = invalidate_refill ? 1'h0 : _GEN_243; // @[TLB.scala 252:34]
  assign _GEN_252 = invalidate_refill ? 1'h0 : _GEN_244; // @[TLB.scala 252:34]
  assign _GEN_253 = _T_1255 ? _GEN_249 : sectored_entries_6_valid_0; // @[TLB.scala 249:72]
  assign _GEN_254 = _T_1255 ? _GEN_250 : sectored_entries_6_valid_1; // @[TLB.scala 249:72]
  assign _GEN_255 = _T_1255 ? _GEN_251 : sectored_entries_6_valid_2; // @[TLB.scala 249:72]
  assign _GEN_256 = _T_1255 ? _GEN_252 : sectored_entries_6_valid_3; // @[TLB.scala 249:72]
  assign _T_1273 = _T_1146 == 3'h7; // @[TLB.scala 249:65]
  assign _GEN_263 = r_sectored_hit ? sectored_entries_7_valid_0 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_264 = r_sectored_hit ? sectored_entries_7_valid_1 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_265 = r_sectored_hit ? sectored_entries_7_valid_2 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_266 = r_sectored_hit ? sectored_entries_7_valid_3 : 1'h0; // @[TLB.scala 250:32]
  assign _GEN_267 = _GEN_995 | _GEN_263; // @[TLB.scala 122:16]
  assign _GEN_268 = _GEN_996 | _GEN_264; // @[TLB.scala 122:16]
  assign _GEN_269 = _GEN_997 | _GEN_265; // @[TLB.scala 122:16]
  assign _GEN_270 = _GEN_998 | _GEN_266; // @[TLB.scala 122:16]
  assign _GEN_275 = invalidate_refill ? 1'h0 : _GEN_267; // @[TLB.scala 252:34]
  assign _GEN_276 = invalidate_refill ? 1'h0 : _GEN_268; // @[TLB.scala 252:34]
  assign _GEN_277 = invalidate_refill ? 1'h0 : _GEN_269; // @[TLB.scala 252:34]
  assign _GEN_278 = invalidate_refill ? 1'h0 : _GEN_270; // @[TLB.scala 252:34]
  assign _GEN_279 = _T_1273 ? _GEN_275 : sectored_entries_7_valid_0; // @[TLB.scala 249:72]
  assign _GEN_280 = _T_1273 ? _GEN_276 : sectored_entries_7_valid_1; // @[TLB.scala 249:72]
  assign _GEN_281 = _T_1273 ? _GEN_277 : sectored_entries_7_valid_2; // @[TLB.scala 249:72]
  assign _GEN_282 = _T_1273 ? _GEN_278 : sectored_entries_7_valid_3; // @[TLB.scala 249:72]
  assign _GEN_291 = _T_1077 ? _GEN_67 : superpage_entries_0_valid_0; // @[TLB.scala 242:54]
  assign _GEN_295 = _T_1077 ? _GEN_71 : superpage_entries_1_valid_0; // @[TLB.scala 242:54]
  assign _GEN_299 = _T_1077 ? _GEN_75 : superpage_entries_2_valid_0; // @[TLB.scala 242:54]
  assign _GEN_303 = _T_1077 ? _GEN_79 : superpage_entries_3_valid_0; // @[TLB.scala 242:54]
  assign _GEN_305 = _T_1077 ? sectored_entries_0_valid_0 : _GEN_97; // @[TLB.scala 242:54]
  assign _GEN_306 = _T_1077 ? sectored_entries_0_valid_1 : _GEN_98; // @[TLB.scala 242:54]
  assign _GEN_307 = _T_1077 ? sectored_entries_0_valid_2 : _GEN_99; // @[TLB.scala 242:54]
  assign _GEN_308 = _T_1077 ? sectored_entries_0_valid_3 : _GEN_100; // @[TLB.scala 242:54]
  assign _GEN_315 = _T_1077 ? sectored_entries_1_valid_0 : _GEN_123; // @[TLB.scala 242:54]
  assign _GEN_316 = _T_1077 ? sectored_entries_1_valid_1 : _GEN_124; // @[TLB.scala 242:54]
  assign _GEN_317 = _T_1077 ? sectored_entries_1_valid_2 : _GEN_125; // @[TLB.scala 242:54]
  assign _GEN_318 = _T_1077 ? sectored_entries_1_valid_3 : _GEN_126; // @[TLB.scala 242:54]
  assign _GEN_325 = _T_1077 ? sectored_entries_2_valid_0 : _GEN_149; // @[TLB.scala 242:54]
  assign _GEN_326 = _T_1077 ? sectored_entries_2_valid_1 : _GEN_150; // @[TLB.scala 242:54]
  assign _GEN_327 = _T_1077 ? sectored_entries_2_valid_2 : _GEN_151; // @[TLB.scala 242:54]
  assign _GEN_328 = _T_1077 ? sectored_entries_2_valid_3 : _GEN_152; // @[TLB.scala 242:54]
  assign _GEN_335 = _T_1077 ? sectored_entries_3_valid_0 : _GEN_175; // @[TLB.scala 242:54]
  assign _GEN_336 = _T_1077 ? sectored_entries_3_valid_1 : _GEN_176; // @[TLB.scala 242:54]
  assign _GEN_337 = _T_1077 ? sectored_entries_3_valid_2 : _GEN_177; // @[TLB.scala 242:54]
  assign _GEN_338 = _T_1077 ? sectored_entries_3_valid_3 : _GEN_178; // @[TLB.scala 242:54]
  assign _GEN_345 = _T_1077 ? sectored_entries_4_valid_0 : _GEN_201; // @[TLB.scala 242:54]
  assign _GEN_346 = _T_1077 ? sectored_entries_4_valid_1 : _GEN_202; // @[TLB.scala 242:54]
  assign _GEN_347 = _T_1077 ? sectored_entries_4_valid_2 : _GEN_203; // @[TLB.scala 242:54]
  assign _GEN_348 = _T_1077 ? sectored_entries_4_valid_3 : _GEN_204; // @[TLB.scala 242:54]
  assign _GEN_355 = _T_1077 ? sectored_entries_5_valid_0 : _GEN_227; // @[TLB.scala 242:54]
  assign _GEN_356 = _T_1077 ? sectored_entries_5_valid_1 : _GEN_228; // @[TLB.scala 242:54]
  assign _GEN_357 = _T_1077 ? sectored_entries_5_valid_2 : _GEN_229; // @[TLB.scala 242:54]
  assign _GEN_358 = _T_1077 ? sectored_entries_5_valid_3 : _GEN_230; // @[TLB.scala 242:54]
  assign _GEN_365 = _T_1077 ? sectored_entries_6_valid_0 : _GEN_253; // @[TLB.scala 242:54]
  assign _GEN_366 = _T_1077 ? sectored_entries_6_valid_1 : _GEN_254; // @[TLB.scala 242:54]
  assign _GEN_367 = _T_1077 ? sectored_entries_6_valid_2 : _GEN_255; // @[TLB.scala 242:54]
  assign _GEN_368 = _T_1077 ? sectored_entries_6_valid_3 : _GEN_256; // @[TLB.scala 242:54]
  assign _GEN_375 = _T_1077 ? sectored_entries_7_valid_0 : _GEN_279; // @[TLB.scala 242:54]
  assign _GEN_376 = _T_1077 ? sectored_entries_7_valid_1 : _GEN_280; // @[TLB.scala 242:54]
  assign _GEN_377 = _T_1077 ? sectored_entries_7_valid_2 : _GEN_281; // @[TLB.scala 242:54]
  assign _GEN_378 = _T_1077 ? sectored_entries_7_valid_3 : _GEN_282; // @[TLB.scala 242:54]
  assign _GEN_387 = io_ptw_resp_bits_homogeneous ? special_entry_valid_0 : _GEN_64; // @[TLB.scala 237:68]
  assign _GEN_391 = io_ptw_resp_bits_homogeneous ? _GEN_291 : superpage_entries_0_valid_0; // @[TLB.scala 237:68]
  assign _GEN_395 = io_ptw_resp_bits_homogeneous ? _GEN_295 : superpage_entries_1_valid_0; // @[TLB.scala 237:68]
  assign _GEN_399 = io_ptw_resp_bits_homogeneous ? _GEN_299 : superpage_entries_2_valid_0; // @[TLB.scala 237:68]
  assign _GEN_403 = io_ptw_resp_bits_homogeneous ? _GEN_303 : superpage_entries_3_valid_0; // @[TLB.scala 237:68]
  assign _GEN_405 = io_ptw_resp_bits_homogeneous ? _GEN_305 : sectored_entries_0_valid_0; // @[TLB.scala 237:68]
  assign _GEN_406 = io_ptw_resp_bits_homogeneous ? _GEN_306 : sectored_entries_0_valid_1; // @[TLB.scala 237:68]
  assign _GEN_407 = io_ptw_resp_bits_homogeneous ? _GEN_307 : sectored_entries_0_valid_2; // @[TLB.scala 237:68]
  assign _GEN_408 = io_ptw_resp_bits_homogeneous ? _GEN_308 : sectored_entries_0_valid_3; // @[TLB.scala 237:68]
  assign _GEN_415 = io_ptw_resp_bits_homogeneous ? _GEN_315 : sectored_entries_1_valid_0; // @[TLB.scala 237:68]
  assign _GEN_416 = io_ptw_resp_bits_homogeneous ? _GEN_316 : sectored_entries_1_valid_1; // @[TLB.scala 237:68]
  assign _GEN_417 = io_ptw_resp_bits_homogeneous ? _GEN_317 : sectored_entries_1_valid_2; // @[TLB.scala 237:68]
  assign _GEN_418 = io_ptw_resp_bits_homogeneous ? _GEN_318 : sectored_entries_1_valid_3; // @[TLB.scala 237:68]
  assign _GEN_425 = io_ptw_resp_bits_homogeneous ? _GEN_325 : sectored_entries_2_valid_0; // @[TLB.scala 237:68]
  assign _GEN_426 = io_ptw_resp_bits_homogeneous ? _GEN_326 : sectored_entries_2_valid_1; // @[TLB.scala 237:68]
  assign _GEN_427 = io_ptw_resp_bits_homogeneous ? _GEN_327 : sectored_entries_2_valid_2; // @[TLB.scala 237:68]
  assign _GEN_428 = io_ptw_resp_bits_homogeneous ? _GEN_328 : sectored_entries_2_valid_3; // @[TLB.scala 237:68]
  assign _GEN_435 = io_ptw_resp_bits_homogeneous ? _GEN_335 : sectored_entries_3_valid_0; // @[TLB.scala 237:68]
  assign _GEN_436 = io_ptw_resp_bits_homogeneous ? _GEN_336 : sectored_entries_3_valid_1; // @[TLB.scala 237:68]
  assign _GEN_437 = io_ptw_resp_bits_homogeneous ? _GEN_337 : sectored_entries_3_valid_2; // @[TLB.scala 237:68]
  assign _GEN_438 = io_ptw_resp_bits_homogeneous ? _GEN_338 : sectored_entries_3_valid_3; // @[TLB.scala 237:68]
  assign _GEN_445 = io_ptw_resp_bits_homogeneous ? _GEN_345 : sectored_entries_4_valid_0; // @[TLB.scala 237:68]
  assign _GEN_446 = io_ptw_resp_bits_homogeneous ? _GEN_346 : sectored_entries_4_valid_1; // @[TLB.scala 237:68]
  assign _GEN_447 = io_ptw_resp_bits_homogeneous ? _GEN_347 : sectored_entries_4_valid_2; // @[TLB.scala 237:68]
  assign _GEN_448 = io_ptw_resp_bits_homogeneous ? _GEN_348 : sectored_entries_4_valid_3; // @[TLB.scala 237:68]
  assign _GEN_455 = io_ptw_resp_bits_homogeneous ? _GEN_355 : sectored_entries_5_valid_0; // @[TLB.scala 237:68]
  assign _GEN_456 = io_ptw_resp_bits_homogeneous ? _GEN_356 : sectored_entries_5_valid_1; // @[TLB.scala 237:68]
  assign _GEN_457 = io_ptw_resp_bits_homogeneous ? _GEN_357 : sectored_entries_5_valid_2; // @[TLB.scala 237:68]
  assign _GEN_458 = io_ptw_resp_bits_homogeneous ? _GEN_358 : sectored_entries_5_valid_3; // @[TLB.scala 237:68]
  assign _GEN_465 = io_ptw_resp_bits_homogeneous ? _GEN_365 : sectored_entries_6_valid_0; // @[TLB.scala 237:68]
  assign _GEN_466 = io_ptw_resp_bits_homogeneous ? _GEN_366 : sectored_entries_6_valid_1; // @[TLB.scala 237:68]
  assign _GEN_467 = io_ptw_resp_bits_homogeneous ? _GEN_367 : sectored_entries_6_valid_2; // @[TLB.scala 237:68]
  assign _GEN_468 = io_ptw_resp_bits_homogeneous ? _GEN_368 : sectored_entries_6_valid_3; // @[TLB.scala 237:68]
  assign _GEN_475 = io_ptw_resp_bits_homogeneous ? _GEN_375 : sectored_entries_7_valid_0; // @[TLB.scala 237:68]
  assign _GEN_476 = io_ptw_resp_bits_homogeneous ? _GEN_376 : sectored_entries_7_valid_1; // @[TLB.scala 237:68]
  assign _GEN_477 = io_ptw_resp_bits_homogeneous ? _GEN_377 : sectored_entries_7_valid_2; // @[TLB.scala 237:68]
  assign _GEN_478 = io_ptw_resp_bits_homogeneous ? _GEN_378 : sectored_entries_7_valid_3; // @[TLB.scala 237:68]
  assign _GEN_487 = io_ptw_resp_valid ? _GEN_387 : special_entry_valid_0; // @[TLB.scala 217:20]
  assign _GEN_491 = io_ptw_resp_valid ? _GEN_391 : superpage_entries_0_valid_0; // @[TLB.scala 217:20]
  assign _GEN_495 = io_ptw_resp_valid ? _GEN_395 : superpage_entries_1_valid_0; // @[TLB.scala 217:20]
  assign _GEN_499 = io_ptw_resp_valid ? _GEN_399 : superpage_entries_2_valid_0; // @[TLB.scala 217:20]
  assign _GEN_503 = io_ptw_resp_valid ? _GEN_403 : superpage_entries_3_valid_0; // @[TLB.scala 217:20]
  assign _GEN_505 = io_ptw_resp_valid ? _GEN_405 : sectored_entries_0_valid_0; // @[TLB.scala 217:20]
  assign _GEN_506 = io_ptw_resp_valid ? _GEN_406 : sectored_entries_0_valid_1; // @[TLB.scala 217:20]
  assign _GEN_507 = io_ptw_resp_valid ? _GEN_407 : sectored_entries_0_valid_2; // @[TLB.scala 217:20]
  assign _GEN_508 = io_ptw_resp_valid ? _GEN_408 : sectored_entries_0_valid_3; // @[TLB.scala 217:20]
  assign _GEN_515 = io_ptw_resp_valid ? _GEN_415 : sectored_entries_1_valid_0; // @[TLB.scala 217:20]
  assign _GEN_516 = io_ptw_resp_valid ? _GEN_416 : sectored_entries_1_valid_1; // @[TLB.scala 217:20]
  assign _GEN_517 = io_ptw_resp_valid ? _GEN_417 : sectored_entries_1_valid_2; // @[TLB.scala 217:20]
  assign _GEN_518 = io_ptw_resp_valid ? _GEN_418 : sectored_entries_1_valid_3; // @[TLB.scala 217:20]
  assign _GEN_525 = io_ptw_resp_valid ? _GEN_425 : sectored_entries_2_valid_0; // @[TLB.scala 217:20]
  assign _GEN_526 = io_ptw_resp_valid ? _GEN_426 : sectored_entries_2_valid_1; // @[TLB.scala 217:20]
  assign _GEN_527 = io_ptw_resp_valid ? _GEN_427 : sectored_entries_2_valid_2; // @[TLB.scala 217:20]
  assign _GEN_528 = io_ptw_resp_valid ? _GEN_428 : sectored_entries_2_valid_3; // @[TLB.scala 217:20]
  assign _GEN_535 = io_ptw_resp_valid ? _GEN_435 : sectored_entries_3_valid_0; // @[TLB.scala 217:20]
  assign _GEN_536 = io_ptw_resp_valid ? _GEN_436 : sectored_entries_3_valid_1; // @[TLB.scala 217:20]
  assign _GEN_537 = io_ptw_resp_valid ? _GEN_437 : sectored_entries_3_valid_2; // @[TLB.scala 217:20]
  assign _GEN_538 = io_ptw_resp_valid ? _GEN_438 : sectored_entries_3_valid_3; // @[TLB.scala 217:20]
  assign _GEN_545 = io_ptw_resp_valid ? _GEN_445 : sectored_entries_4_valid_0; // @[TLB.scala 217:20]
  assign _GEN_546 = io_ptw_resp_valid ? _GEN_446 : sectored_entries_4_valid_1; // @[TLB.scala 217:20]
  assign _GEN_547 = io_ptw_resp_valid ? _GEN_447 : sectored_entries_4_valid_2; // @[TLB.scala 217:20]
  assign _GEN_548 = io_ptw_resp_valid ? _GEN_448 : sectored_entries_4_valid_3; // @[TLB.scala 217:20]
  assign _GEN_555 = io_ptw_resp_valid ? _GEN_455 : sectored_entries_5_valid_0; // @[TLB.scala 217:20]
  assign _GEN_556 = io_ptw_resp_valid ? _GEN_456 : sectored_entries_5_valid_1; // @[TLB.scala 217:20]
  assign _GEN_557 = io_ptw_resp_valid ? _GEN_457 : sectored_entries_5_valid_2; // @[TLB.scala 217:20]
  assign _GEN_558 = io_ptw_resp_valid ? _GEN_458 : sectored_entries_5_valid_3; // @[TLB.scala 217:20]
  assign _GEN_565 = io_ptw_resp_valid ? _GEN_465 : sectored_entries_6_valid_0; // @[TLB.scala 217:20]
  assign _GEN_566 = io_ptw_resp_valid ? _GEN_466 : sectored_entries_6_valid_1; // @[TLB.scala 217:20]
  assign _GEN_567 = io_ptw_resp_valid ? _GEN_467 : sectored_entries_6_valid_2; // @[TLB.scala 217:20]
  assign _GEN_568 = io_ptw_resp_valid ? _GEN_468 : sectored_entries_6_valid_3; // @[TLB.scala 217:20]
  assign _GEN_575 = io_ptw_resp_valid ? _GEN_475 : sectored_entries_7_valid_0; // @[TLB.scala 217:20]
  assign _GEN_576 = io_ptw_resp_valid ? _GEN_476 : sectored_entries_7_valid_1; // @[TLB.scala 217:20]
  assign _GEN_577 = io_ptw_resp_valid ? _GEN_477 : sectored_entries_7_valid_2; // @[TLB.scala 217:20]
  assign _GEN_578 = io_ptw_resp_valid ? _GEN_478 : sectored_entries_7_valid_3; // @[TLB.scala 217:20]
  assign _T_1761 = {OptimizationBarrier_19_io_y_ae,OptimizationBarrier_18_io_y_ae,OptimizationBarrier_17_io_y_ae,OptimizationBarrier_16_io_y_ae,OptimizationBarrier_15_io_y_ae,OptimizationBarrier_14_io_y_ae}; // @[Cat.scala 29:58]
  assign ptw_ae_array = {1'h0,OptimizationBarrier_26_io_y_ae,OptimizationBarrier_25_io_y_ae,OptimizationBarrier_24_io_y_ae,OptimizationBarrier_23_io_y_ae,OptimizationBarrier_22_io_y_ae,OptimizationBarrier_21_io_y_ae,OptimizationBarrier_20_io_y_ae,_T_1761}; // @[Cat.scala 29:58]
  assign _T_1775 = {OptimizationBarrier_19_io_y_u,OptimizationBarrier_18_io_y_u,OptimizationBarrier_17_io_y_u,OptimizationBarrier_16_io_y_u,OptimizationBarrier_15_io_y_u,OptimizationBarrier_14_io_y_u}; // @[Cat.scala 29:58]
  assign _T_1782 = {OptimizationBarrier_26_io_y_u,OptimizationBarrier_25_io_y_u,OptimizationBarrier_24_io_y_u,OptimizationBarrier_23_io_y_u,OptimizationBarrier_22_io_y_u,OptimizationBarrier_21_io_y_u,OptimizationBarrier_20_io_y_u,_T_1775}; // @[Cat.scala 29:58]
  assign priv_x_ok = priv_s ? ~_T_1782 : _T_1782; // @[TLB.scala 262:22]
  assign _T_1839 = {OptimizationBarrier_19_io_y_sx,OptimizationBarrier_18_io_y_sx,OptimizationBarrier_17_io_y_sx,OptimizationBarrier_16_io_y_sx,OptimizationBarrier_15_io_y_sx,OptimizationBarrier_14_io_y_sx}; // @[Cat.scala 29:58]
  assign _T_1846 = {OptimizationBarrier_26_io_y_sx,OptimizationBarrier_25_io_y_sx,OptimizationBarrier_24_io_y_sx,OptimizationBarrier_23_io_y_sx,OptimizationBarrier_22_io_y_sx,OptimizationBarrier_21_io_y_sx,OptimizationBarrier_20_io_y_sx,_T_1839}; // @[Cat.scala 29:58]
  assign _T_1875 = priv_x_ok & _T_1846; // @[TLB.scala 265:39]
  assign x_array = {1'h1,_T_1875}; // @[Cat.scala 29:58]
  assign _T_1907 = prot_x ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_1912 = {OptimizationBarrier_32_io_y_px,OptimizationBarrier_31_io_y_px,OptimizationBarrier_30_io_y_px,OptimizationBarrier_29_io_y_px,OptimizationBarrier_28_io_y_px,OptimizationBarrier_27_io_y_px}; // @[Cat.scala 29:58]
  assign _T_1919 = {_T_1907,OptimizationBarrier_38_io_y_px,OptimizationBarrier_37_io_y_px,OptimizationBarrier_36_io_y_px,OptimizationBarrier_35_io_y_px,OptimizationBarrier_34_io_y_px,OptimizationBarrier_33_io_y_px,_T_1912}; // @[Cat.scala 29:58]
  assign px_array = _T_1919 & ~ptw_ae_array; // @[TLB.scala 268:87]
  assign _T_1935 = cacheable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_1940 = {OptimizationBarrier_32_io_y_c,OptimizationBarrier_31_io_y_c,OptimizationBarrier_30_io_y_c,OptimizationBarrier_29_io_y_c,OptimizationBarrier_28_io_y_c,OptimizationBarrier_27_io_y_c}; // @[Cat.scala 29:58]
  assign c_array = {_T_1935,OptimizationBarrier_38_io_y_c,OptimizationBarrier_37_io_y_c,OptimizationBarrier_36_io_y_c,OptimizationBarrier_35_io_y_c,OptimizationBarrier_34_io_y_c,OptimizationBarrier_33_io_y_c,_T_1940}; // @[Cat.scala 29:58]
  assign _T_2005 = io_req_bits_vaddr & 40'hc000000000; // @[TLB.scala 285:43]
  assign _T_2007 = _T_2005 == 40'h0; // @[TLB.scala 286:61]
  assign _T_2008 = _T_2005 == 40'hc000000000; // @[TLB.scala 286:82]
  assign _T_2009 = _T_2007 | _T_2008; // @[TLB.scala 286:67]
  assign bad_va = vm_enabled & ~_T_2009; // @[TLB.scala 280:117]
  assign _T_2112 = x_array | ptw_ae_array; // @[TLB.scala 318:33]
  assign pf_inst_array = ~_T_2112; // @[TLB.scala 318:23]
  assign tlb_hit = |real_hits; // @[TLB.scala 320:27]
  assign _T_2114 = vm_enabled & ~bad_va; // @[TLB.scala 321:29]
  assign tlb_miss = _T_2114 & ~tlb_hit; // @[TLB.scala 321:40]
  assign _T_2118 = io_req_valid & vm_enabled; // @[TLB.scala 325:22]
  assign _T_2119 = sector_hits_0 | sector_hits_1; // @[package.scala 64:59]
  assign _T_2120 = _T_2119 | sector_hits_2; // @[package.scala 64:59]
  assign _T_2121 = _T_2120 | sector_hits_3; // @[package.scala 64:59]
  assign _T_2122 = _T_2121 | sector_hits_4; // @[package.scala 64:59]
  assign _T_2123 = _T_2122 | sector_hits_5; // @[package.scala 64:59]
  assign _T_2124 = _T_2123 | sector_hits_6; // @[package.scala 64:59]
  assign _T_2125 = _T_2124 | sector_hits_7; // @[package.scala 64:59]
  assign _T_2132 = {sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0}; // @[Cat.scala 29:58]
  assign _T_2135 = |_T_2132[7:4]; // @[OneHot.scala 32:14]
  assign _T_2136 = _T_2132[7:4] | _T_2132[3:0]; // @[OneHot.scala 32:28]
  assign _T_2139 = |_T_2136[3:2]; // @[OneHot.scala 32:14]
  assign _T_2140 = _T_2136[3:2] | _T_2136[1:0]; // @[OneHot.scala 32:28]
  assign _T_2143 = {_T_2135,_T_2139,_T_2140[1]}; // @[Cat.scala 29:58]
  assign _T_2157 = _T_2143[1] ? ~_T_2143[0] : _T_2116[4]; // @[Replacement.scala 193:16]
  assign _T_2161 = _T_2143[1] ? _T_2116[3] : ~_T_2143[0]; // @[Replacement.scala 196:16]
  assign _T_2163 = {~_T_2143[1],_T_2157,_T_2161}; // @[Cat.scala 29:58]
  assign _T_2164 = _T_2143[2] ? _T_2163 : _T_2116[5:3]; // @[Replacement.scala 193:16]
  assign _T_2173 = _T_2143[1] ? ~_T_2143[0] : _T_2116[1]; // @[Replacement.scala 193:16]
  assign _T_2177 = _T_2143[1] ? _T_2116[0] : ~_T_2143[0]; // @[Replacement.scala 196:16]
  assign _T_2179 = {~_T_2143[1],_T_2173,_T_2177}; // @[Cat.scala 29:58]
  assign _T_2180 = _T_2143[2] ? _T_2116[2:0] : _T_2179; // @[Replacement.scala 196:16]
  assign _T_2182 = {~_T_2143[2],_T_2164,_T_2180}; // @[Cat.scala 29:58]
  assign _T_2183 = superpage_hits_0 | superpage_hits_1; // @[package.scala 64:59]
  assign _T_2184 = _T_2183 | superpage_hits_2; // @[package.scala 64:59]
  assign _T_2185 = _T_2184 | superpage_hits_3; // @[package.scala 64:59]
  assign _T_2188 = {superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; // @[Cat.scala 29:58]
  assign _T_2191 = |_T_2188[3:2]; // @[OneHot.scala 32:14]
  assign _T_2192 = _T_2188[3:2] | _T_2188[1:0]; // @[OneHot.scala 32:28]
  assign _T_2194 = {_T_2191,_T_2192[1]}; // @[Cat.scala 29:58]
  assign _T_2203 = _T_2194[1] ? ~_T_2194[0] : _T_2117[1]; // @[Replacement.scala 193:16]
  assign _T_2207 = _T_2194[1] ? _T_2117[0] : ~_T_2194[0]; // @[Replacement.scala 196:16]
  assign _T_2209 = {~_T_2194[1],_T_2203,_T_2207}; // @[Cat.scala 29:58]
  assign _T_2219 = real_hits[1] | real_hits[2]; // @[Misc.scala 182:16]
  assign _T_2221 = real_hits[1] & real_hits[2]; // @[Misc.scala 182:61]
  assign _T_2223 = real_hits[0] | _T_2219; // @[Misc.scala 182:16]
  assign _T_2225 = real_hits[0] & _T_2219; // @[Misc.scala 182:61]
  assign _T_2226 = _T_2221 | _T_2225; // @[Misc.scala 182:49]
  assign _T_2235 = real_hits[4] | real_hits[5]; // @[Misc.scala 182:16]
  assign _T_2237 = real_hits[4] & real_hits[5]; // @[Misc.scala 182:61]
  assign _T_2239 = real_hits[3] | _T_2235; // @[Misc.scala 182:16]
  assign _T_2241 = real_hits[3] & _T_2235; // @[Misc.scala 182:61]
  assign _T_2242 = _T_2237 | _T_2241; // @[Misc.scala 182:49]
  assign _T_2243 = _T_2223 | _T_2239; // @[Misc.scala 182:16]
  assign _T_2244 = _T_2226 | _T_2242; // @[Misc.scala 182:37]
  assign _T_2245 = _T_2223 & _T_2239; // @[Misc.scala 182:61]
  assign _T_2246 = _T_2244 | _T_2245; // @[Misc.scala 182:49]
  assign _T_2256 = real_hits[7] | real_hits[8]; // @[Misc.scala 182:16]
  assign _T_2258 = real_hits[7] & real_hits[8]; // @[Misc.scala 182:61]
  assign _T_2260 = real_hits[6] | _T_2256; // @[Misc.scala 182:16]
  assign _T_2262 = real_hits[6] & _T_2256; // @[Misc.scala 182:61]
  assign _T_2263 = _T_2258 | _T_2262; // @[Misc.scala 182:49]
  assign _T_2270 = real_hits[9] | real_hits[10]; // @[Misc.scala 182:16]
  assign _T_2272 = real_hits[9] & real_hits[10]; // @[Misc.scala 182:61]
  assign _T_2279 = real_hits[11] | real_hits[12]; // @[Misc.scala 182:16]
  assign _T_2281 = real_hits[11] & real_hits[12]; // @[Misc.scala 182:61]
  assign _T_2283 = _T_2270 | _T_2279; // @[Misc.scala 182:16]
  assign _T_2284 = _T_2272 | _T_2281; // @[Misc.scala 182:37]
  assign _T_2285 = _T_2270 & _T_2279; // @[Misc.scala 182:61]
  assign _T_2286 = _T_2284 | _T_2285; // @[Misc.scala 182:49]
  assign _T_2287 = _T_2260 | _T_2283; // @[Misc.scala 182:16]
  assign _T_2288 = _T_2263 | _T_2286; // @[Misc.scala 182:37]
  assign _T_2289 = _T_2260 & _T_2283; // @[Misc.scala 182:61]
  assign _T_2290 = _T_2288 | _T_2289; // @[Misc.scala 182:49]
  assign _T_2292 = _T_2246 | _T_2290; // @[Misc.scala 182:37]
  assign _T_2293 = _T_2243 & _T_2287; // @[Misc.scala 182:61]
  assign multipleHits = _T_2292 | _T_2293; // @[Misc.scala 182:49]
  assign _T_2303 = pf_inst_array & hits; // @[TLB.scala 340:47]
  assign _T_2304 = |_T_2303; // @[TLB.scala 340:55]
  assign _T_2311 = ~px_array & hits; // @[TLB.scala 343:33]
  assign _T_2317 = c_array & hits; // @[TLB.scala 347:33]
  assign _T_2324 = io_ptw_resp_valid | tlb_miss; // @[TLB.scala 350:29]
  assign _T_2330 = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37]
  assign _T_2331 = _T_2330 & tlb_miss; // @[TLB.scala 359:25]
  assign _T_2337 = _T_2117[2] ? _T_2117[1] : _T_2117[0]; // @[Replacement.scala 240:16]
  assign _T_2338 = {_T_2117[2],_T_2337}; // @[Cat.scala 29:58]
  assign _T_2341 = {superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[Cat.scala 29:58]
  assign _T_2342 = &_T_2341; // @[TLB.scala 407:16]
  assign _T_2344 = ~_T_2341[0]; // @[OneHot.scala 47:40]
  assign _T_2345 = ~_T_2341[1]; // @[OneHot.scala 47:40]
  assign _T_2346 = ~_T_2341[2]; // @[OneHot.scala 47:40]
  assign _T_2360 = _T_2116[5] ? _T_2116[4] : _T_2116[3]; // @[Replacement.scala 240:16]
  assign _T_2361 = {_T_2116[5],_T_2360}; // @[Cat.scala 29:58]
  assign _T_2367 = _T_2116[2] ? _T_2116[1] : _T_2116[0]; // @[Replacement.scala 240:16]
  assign _T_2368 = {_T_2116[2],_T_2367}; // @[Cat.scala 29:58]
  assign _T_2369 = _T_2116[6] ? _T_2361 : _T_2368; // @[Replacement.scala 240:16]
  assign _T_2370 = {_T_2116[6],_T_2369}; // @[Cat.scala 29:58]
  assign _T_2401 = {_T_461,_T_455,_T_449,_T_443,_T_437,_T_431,_T_425,_T_419}; // @[Cat.scala 29:58]
  assign _T_2402 = &_T_2401; // @[TLB.scala 407:16]
  assign _T_2404 = ~_T_2401[0]; // @[OneHot.scala 47:40]
  assign _T_2405 = ~_T_2401[1]; // @[OneHot.scala 47:40]
  assign _T_2406 = ~_T_2401[2]; // @[OneHot.scala 47:40]
  assign _T_2407 = ~_T_2401[3]; // @[OneHot.scala 47:40]
  assign _T_2408 = ~_T_2401[4]; // @[OneHot.scala 47:40]
  assign _T_2409 = ~_T_2401[5]; // @[OneHot.scala 47:40]
  assign _T_2410 = ~_T_2401[6]; // @[OneHot.scala 47:40]
  assign _T_2447 = state == 2'h2; // @[TLB.scala 373:17]
  assign _T_2448 = _T_2447 & io_sfence_valid; // @[TLB.scala 373:28]
  assign _T_2451 = io_sfence_bits_addr[38:12] == vpn; // @[TLB.scala 381:72]
  assign _T_2452 = ~io_sfence_bits_rs1 | _T_2451; // @[TLB.scala 381:34]
  assign _T_2454 = _T_2452 | reset; // @[TLB.scala 381:13]
  assign _T_2462 = _T_420[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_681 = sectored_entries_0_data_0[13] ? _GEN_505 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_682 = sectored_entries_0_data_1[13] ? _GEN_506 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_683 = sectored_entries_0_data_2[13] ? _GEN_507 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_684 = sectored_entries_0_data_3[13] ? _GEN_508 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_685 = io_sfence_bits_rs2 & _GEN_681; // @[TLB.scala 384:40]
  assign _GEN_686 = io_sfence_bits_rs2 & _GEN_682; // @[TLB.scala 384:40]
  assign _GEN_687 = io_sfence_bits_rs2 & _GEN_683; // @[TLB.scala 384:40]
  assign _GEN_688 = io_sfence_bits_rs2 & _GEN_684; // @[TLB.scala 384:40]
  assign _T_2617 = _T_426[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_709 = sectored_entries_1_data_0[13] ? _GEN_515 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_710 = sectored_entries_1_data_1[13] ? _GEN_516 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_711 = sectored_entries_1_data_2[13] ? _GEN_517 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_712 = sectored_entries_1_data_3[13] ? _GEN_518 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_713 = io_sfence_bits_rs2 & _GEN_709; // @[TLB.scala 384:40]
  assign _GEN_714 = io_sfence_bits_rs2 & _GEN_710; // @[TLB.scala 384:40]
  assign _GEN_715 = io_sfence_bits_rs2 & _GEN_711; // @[TLB.scala 384:40]
  assign _GEN_716 = io_sfence_bits_rs2 & _GEN_712; // @[TLB.scala 384:40]
  assign _T_2772 = _T_432[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_737 = sectored_entries_2_data_0[13] ? _GEN_525 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_738 = sectored_entries_2_data_1[13] ? _GEN_526 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_739 = sectored_entries_2_data_2[13] ? _GEN_527 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_740 = sectored_entries_2_data_3[13] ? _GEN_528 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_741 = io_sfence_bits_rs2 & _GEN_737; // @[TLB.scala 384:40]
  assign _GEN_742 = io_sfence_bits_rs2 & _GEN_738; // @[TLB.scala 384:40]
  assign _GEN_743 = io_sfence_bits_rs2 & _GEN_739; // @[TLB.scala 384:40]
  assign _GEN_744 = io_sfence_bits_rs2 & _GEN_740; // @[TLB.scala 384:40]
  assign _T_2927 = _T_438[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_765 = sectored_entries_3_data_0[13] ? _GEN_535 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_766 = sectored_entries_3_data_1[13] ? _GEN_536 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_767 = sectored_entries_3_data_2[13] ? _GEN_537 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_768 = sectored_entries_3_data_3[13] ? _GEN_538 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_769 = io_sfence_bits_rs2 & _GEN_765; // @[TLB.scala 384:40]
  assign _GEN_770 = io_sfence_bits_rs2 & _GEN_766; // @[TLB.scala 384:40]
  assign _GEN_771 = io_sfence_bits_rs2 & _GEN_767; // @[TLB.scala 384:40]
  assign _GEN_772 = io_sfence_bits_rs2 & _GEN_768; // @[TLB.scala 384:40]
  assign _T_3082 = _T_444[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_793 = sectored_entries_4_data_0[13] ? _GEN_545 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_794 = sectored_entries_4_data_1[13] ? _GEN_546 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_795 = sectored_entries_4_data_2[13] ? _GEN_547 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_796 = sectored_entries_4_data_3[13] ? _GEN_548 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_797 = io_sfence_bits_rs2 & _GEN_793; // @[TLB.scala 384:40]
  assign _GEN_798 = io_sfence_bits_rs2 & _GEN_794; // @[TLB.scala 384:40]
  assign _GEN_799 = io_sfence_bits_rs2 & _GEN_795; // @[TLB.scala 384:40]
  assign _GEN_800 = io_sfence_bits_rs2 & _GEN_796; // @[TLB.scala 384:40]
  assign _T_3237 = _T_450[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_821 = sectored_entries_5_data_0[13] ? _GEN_555 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_822 = sectored_entries_5_data_1[13] ? _GEN_556 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_823 = sectored_entries_5_data_2[13] ? _GEN_557 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_824 = sectored_entries_5_data_3[13] ? _GEN_558 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_825 = io_sfence_bits_rs2 & _GEN_821; // @[TLB.scala 384:40]
  assign _GEN_826 = io_sfence_bits_rs2 & _GEN_822; // @[TLB.scala 384:40]
  assign _GEN_827 = io_sfence_bits_rs2 & _GEN_823; // @[TLB.scala 384:40]
  assign _GEN_828 = io_sfence_bits_rs2 & _GEN_824; // @[TLB.scala 384:40]
  assign _T_3392 = _T_456[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_849 = sectored_entries_6_data_0[13] ? _GEN_565 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_850 = sectored_entries_6_data_1[13] ? _GEN_566 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_851 = sectored_entries_6_data_2[13] ? _GEN_567 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_852 = sectored_entries_6_data_3[13] ? _GEN_568 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_853 = io_sfence_bits_rs2 & _GEN_849; // @[TLB.scala 384:40]
  assign _GEN_854 = io_sfence_bits_rs2 & _GEN_850; // @[TLB.scala 384:40]
  assign _GEN_855 = io_sfence_bits_rs2 & _GEN_851; // @[TLB.scala 384:40]
  assign _GEN_856 = io_sfence_bits_rs2 & _GEN_852; // @[TLB.scala 384:40]
  assign _T_3547 = _T_462[26:18] == 9'h0; // @[TLB.scala 135:61]
  assign _GEN_877 = sectored_entries_7_data_0[13] ? _GEN_575 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_878 = sectored_entries_7_data_1[13] ? _GEN_576 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_879 = sectored_entries_7_data_2[13] ? _GEN_577 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_880 = sectored_entries_7_data_3[13] ? _GEN_578 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_881 = io_sfence_bits_rs2 & _GEN_877; // @[TLB.scala 384:40]
  assign _GEN_882 = io_sfence_bits_rs2 & _GEN_878; // @[TLB.scala 384:40]
  assign _GEN_883 = io_sfence_bits_rs2 & _GEN_879; // @[TLB.scala 384:40]
  assign _GEN_884 = io_sfence_bits_rs2 & _GEN_880; // @[TLB.scala 384:40]
  assign _GEN_890 = superpage_entries_0_data_0[13] ? _GEN_491 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_891 = io_sfence_bits_rs2 & _GEN_890; // @[TLB.scala 384:40]
  assign _GEN_894 = superpage_entries_1_data_0[13] ? _GEN_495 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_895 = io_sfence_bits_rs2 & _GEN_894; // @[TLB.scala 384:40]
  assign _GEN_898 = superpage_entries_2_data_0[13] ? _GEN_499 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_899 = io_sfence_bits_rs2 & _GEN_898; // @[TLB.scala 384:40]
  assign _GEN_902 = superpage_entries_3_data_0[13] ? _GEN_503 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_903 = io_sfence_bits_rs2 & _GEN_902; // @[TLB.scala 384:40]
  assign _GEN_906 = special_entry_data_0[13] ? _GEN_487 : 1'h0; // @[TLB.scala 143:19]
  assign _GEN_907 = io_sfence_bits_rs2 & _GEN_906; // @[TLB.scala 384:40]
  assign _T_3897 = multipleHits | reset; // @[TLB.scala 388:24]
  assign io_req_ready = state == 2'h0; // @[TLB.scala 337:16]
  assign io_resp_miss = _T_2324 | multipleHits; // @[TLB.scala 350:16]
  assign io_resp_paddr = {ppn,io_req_bits_vaddr[11:0]}; // @[TLB.scala 351:17]
  assign io_resp_pf_inst = bad_va | _T_2304; // @[TLB.scala 340:19]
  assign io_resp_ae_inst = |_T_2311; // @[TLB.scala 343:19]
  assign io_resp_cacheable = |_T_2317; // @[TLB.scala 347:21]
  assign io_ptw_req_valid = state == 2'h1; // @[TLB.scala 353:20]
  assign io_ptw_req_bits_valid = ~io_kill; // @[TLB.scala 354:25]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[TLB.scala 355:29]
  assign OptimizationBarrier_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_u = special_entry_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_ae = special_entry_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_sw = special_entry_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_sx = special_entry_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_sr = special_entry_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_pw = special_entry_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_px = special_entry_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_pr = special_entry_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_ppp = special_entry_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_pal = special_entry_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_paa = special_entry_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_eff = special_entry_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_io_x_c = special_entry_data_0[1]; // @[package.scala 244:18]
  assign pmp_io_prv = mpu_priv[1:0]; // @[TLB.scala 194:14]
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask; // @[TLB.scala 193:14]
  assign pmp_io_addr = mpu_physaddr[31:0]; // @[TLB.scala 191:15]
  assign OptimizationBarrier_1_io_x_ppn = _GEN_35[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_u = _GEN_35[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_ae = _GEN_35[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_sw = _GEN_35[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_sx = _GEN_35[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_sr = _GEN_35[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_pw = _GEN_35[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_px = _GEN_35[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_pr = _GEN_35[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_ppp = _GEN_35[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_pal = _GEN_35[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_paa = _GEN_35[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_eff = _GEN_35[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_1_io_x_c = _GEN_35[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_ppn = _GEN_39[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_u = _GEN_39[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_ae = _GEN_39[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_sw = _GEN_39[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_sx = _GEN_39[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_sr = _GEN_39[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_pw = _GEN_39[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_px = _GEN_39[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_pr = _GEN_39[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_ppp = _GEN_39[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_pal = _GEN_39[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_paa = _GEN_39[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_eff = _GEN_39[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_2_io_x_c = _GEN_39[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_ppn = _GEN_43[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_u = _GEN_43[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_ae = _GEN_43[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_sw = _GEN_43[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_sx = _GEN_43[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_sr = _GEN_43[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_pw = _GEN_43[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_px = _GEN_43[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_pr = _GEN_43[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_ppp = _GEN_43[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_pal = _GEN_43[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_paa = _GEN_43[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_eff = _GEN_43[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_3_io_x_c = _GEN_43[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_ppn = _GEN_47[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_u = _GEN_47[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_ae = _GEN_47[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_sw = _GEN_47[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_sx = _GEN_47[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_sr = _GEN_47[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_pw = _GEN_47[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_px = _GEN_47[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_pr = _GEN_47[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_ppp = _GEN_47[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_pal = _GEN_47[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_paa = _GEN_47[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_eff = _GEN_47[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_4_io_x_c = _GEN_47[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_ppn = _GEN_51[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_u = _GEN_51[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_ae = _GEN_51[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_sw = _GEN_51[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_sx = _GEN_51[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_sr = _GEN_51[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_pw = _GEN_51[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_px = _GEN_51[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_pr = _GEN_51[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_ppp = _GEN_51[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_pal = _GEN_51[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_paa = _GEN_51[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_eff = _GEN_51[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_5_io_x_c = _GEN_51[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_ppn = _GEN_55[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_u = _GEN_55[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_ae = _GEN_55[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_sw = _GEN_55[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_sx = _GEN_55[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_sr = _GEN_55[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_pw = _GEN_55[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_px = _GEN_55[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_pr = _GEN_55[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_ppp = _GEN_55[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_pal = _GEN_55[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_paa = _GEN_55[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_eff = _GEN_55[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_6_io_x_c = _GEN_55[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_ppn = _GEN_59[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_u = _GEN_59[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_ae = _GEN_59[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_sw = _GEN_59[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_sx = _GEN_59[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_sr = _GEN_59[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_pw = _GEN_59[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_px = _GEN_59[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_pr = _GEN_59[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_ppp = _GEN_59[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_pal = _GEN_59[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_paa = _GEN_59[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_eff = _GEN_59[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_7_io_x_c = _GEN_59[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_ppn = _GEN_63[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_u = _GEN_63[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_ae = _GEN_63[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_sw = _GEN_63[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_sx = _GEN_63[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_sr = _GEN_63[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_pw = _GEN_63[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_px = _GEN_63[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_pr = _GEN_63[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_ppp = _GEN_63[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_pal = _GEN_63[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_paa = _GEN_63[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_eff = _GEN_63[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_8_io_x_c = _GEN_63[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_u = superpage_entries_0_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_ae = superpage_entries_0_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_sw = superpage_entries_0_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_sx = superpage_entries_0_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_sr = superpage_entries_0_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_pw = superpage_entries_0_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_px = superpage_entries_0_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_pr = superpage_entries_0_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_ppp = superpage_entries_0_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_9_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_u = superpage_entries_1_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_ae = superpage_entries_1_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_sw = superpage_entries_1_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_sx = superpage_entries_1_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_sr = superpage_entries_1_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_pw = superpage_entries_1_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_px = superpage_entries_1_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_pr = superpage_entries_1_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_ppp = superpage_entries_1_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_10_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_u = superpage_entries_2_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_ae = superpage_entries_2_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_sw = superpage_entries_2_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_sx = superpage_entries_2_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_sr = superpage_entries_2_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_pw = superpage_entries_2_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_px = superpage_entries_2_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_pr = superpage_entries_2_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_ppp = superpage_entries_2_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_11_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_u = superpage_entries_3_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_ae = superpage_entries_3_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_sw = superpage_entries_3_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_sx = superpage_entries_3_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_sr = superpage_entries_3_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_pw = superpage_entries_3_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_px = superpage_entries_3_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_pr = superpage_entries_3_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_ppp = superpage_entries_3_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_12_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_u = special_entry_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_ae = special_entry_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_sw = special_entry_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_sx = special_entry_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_sr = special_entry_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_pw = special_entry_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_px = special_entry_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_pr = special_entry_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_ppp = special_entry_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_pal = special_entry_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_paa = special_entry_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_eff = special_entry_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_13_io_x_c = special_entry_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_ppn = _GEN_35[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_u = _GEN_35[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_ae = _GEN_35[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_sw = _GEN_35[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_sx = _GEN_35[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_sr = _GEN_35[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_pw = _GEN_35[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_px = _GEN_35[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_pr = _GEN_35[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_ppp = _GEN_35[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_pal = _GEN_35[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_paa = _GEN_35[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_eff = _GEN_35[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_14_io_x_c = _GEN_35[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_ppn = _GEN_39[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_u = _GEN_39[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_ae = _GEN_39[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_sw = _GEN_39[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_sx = _GEN_39[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_sr = _GEN_39[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_pw = _GEN_39[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_px = _GEN_39[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_pr = _GEN_39[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_ppp = _GEN_39[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_pal = _GEN_39[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_paa = _GEN_39[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_eff = _GEN_39[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_15_io_x_c = _GEN_39[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_ppn = _GEN_43[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_u = _GEN_43[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_ae = _GEN_43[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_sw = _GEN_43[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_sx = _GEN_43[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_sr = _GEN_43[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_pw = _GEN_43[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_px = _GEN_43[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_pr = _GEN_43[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_ppp = _GEN_43[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_pal = _GEN_43[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_paa = _GEN_43[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_eff = _GEN_43[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_16_io_x_c = _GEN_43[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_ppn = _GEN_47[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_u = _GEN_47[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_ae = _GEN_47[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_sw = _GEN_47[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_sx = _GEN_47[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_sr = _GEN_47[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_pw = _GEN_47[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_px = _GEN_47[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_pr = _GEN_47[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_ppp = _GEN_47[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_pal = _GEN_47[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_paa = _GEN_47[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_eff = _GEN_47[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_17_io_x_c = _GEN_47[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_ppn = _GEN_51[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_u = _GEN_51[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_ae = _GEN_51[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_sw = _GEN_51[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_sx = _GEN_51[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_sr = _GEN_51[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_pw = _GEN_51[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_px = _GEN_51[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_pr = _GEN_51[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_ppp = _GEN_51[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_pal = _GEN_51[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_paa = _GEN_51[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_eff = _GEN_51[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_18_io_x_c = _GEN_51[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_ppn = _GEN_55[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_u = _GEN_55[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_ae = _GEN_55[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_sw = _GEN_55[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_sx = _GEN_55[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_sr = _GEN_55[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_pw = _GEN_55[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_px = _GEN_55[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_pr = _GEN_55[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_ppp = _GEN_55[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_pal = _GEN_55[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_paa = _GEN_55[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_eff = _GEN_55[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_19_io_x_c = _GEN_55[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_ppn = _GEN_59[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_u = _GEN_59[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_ae = _GEN_59[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_sw = _GEN_59[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_sx = _GEN_59[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_sr = _GEN_59[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_pw = _GEN_59[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_px = _GEN_59[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_pr = _GEN_59[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_ppp = _GEN_59[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_pal = _GEN_59[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_paa = _GEN_59[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_eff = _GEN_59[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_20_io_x_c = _GEN_59[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_ppn = _GEN_63[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_u = _GEN_63[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_ae = _GEN_63[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_sw = _GEN_63[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_sx = _GEN_63[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_sr = _GEN_63[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_pw = _GEN_63[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_px = _GEN_63[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_pr = _GEN_63[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_ppp = _GEN_63[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_pal = _GEN_63[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_paa = _GEN_63[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_eff = _GEN_63[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_21_io_x_c = _GEN_63[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_u = superpage_entries_0_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_ae = superpage_entries_0_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_sw = superpage_entries_0_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_sx = superpage_entries_0_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_sr = superpage_entries_0_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_pw = superpage_entries_0_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_px = superpage_entries_0_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_pr = superpage_entries_0_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_ppp = superpage_entries_0_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_22_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_u = superpage_entries_1_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_ae = superpage_entries_1_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_sw = superpage_entries_1_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_sx = superpage_entries_1_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_sr = superpage_entries_1_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_pw = superpage_entries_1_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_px = superpage_entries_1_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_pr = superpage_entries_1_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_ppp = superpage_entries_1_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_23_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_u = superpage_entries_2_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_ae = superpage_entries_2_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_sw = superpage_entries_2_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_sx = superpage_entries_2_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_sr = superpage_entries_2_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_pw = superpage_entries_2_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_px = superpage_entries_2_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_pr = superpage_entries_2_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_ppp = superpage_entries_2_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_24_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_u = superpage_entries_3_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_ae = superpage_entries_3_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_sw = superpage_entries_3_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_sx = superpage_entries_3_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_sr = superpage_entries_3_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_pw = superpage_entries_3_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_px = superpage_entries_3_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_pr = superpage_entries_3_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_ppp = superpage_entries_3_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_25_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_u = special_entry_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_ae = special_entry_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_sw = special_entry_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_sx = special_entry_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_sr = special_entry_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_pw = special_entry_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_px = special_entry_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_pr = special_entry_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_ppp = special_entry_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_pal = special_entry_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_paa = special_entry_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_eff = special_entry_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_26_io_x_c = special_entry_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_ppn = _GEN_35[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_u = _GEN_35[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_ae = _GEN_35[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_sw = _GEN_35[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_sx = _GEN_35[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_sr = _GEN_35[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_pw = _GEN_35[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_px = _GEN_35[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_pr = _GEN_35[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_ppp = _GEN_35[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_pal = _GEN_35[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_paa = _GEN_35[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_eff = _GEN_35[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_27_io_x_c = _GEN_35[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_ppn = _GEN_39[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_u = _GEN_39[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_ae = _GEN_39[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_sw = _GEN_39[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_sx = _GEN_39[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_sr = _GEN_39[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_pw = _GEN_39[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_px = _GEN_39[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_pr = _GEN_39[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_ppp = _GEN_39[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_pal = _GEN_39[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_paa = _GEN_39[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_eff = _GEN_39[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_28_io_x_c = _GEN_39[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_ppn = _GEN_43[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_u = _GEN_43[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_ae = _GEN_43[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_sw = _GEN_43[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_sx = _GEN_43[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_sr = _GEN_43[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_pw = _GEN_43[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_px = _GEN_43[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_pr = _GEN_43[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_ppp = _GEN_43[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_pal = _GEN_43[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_paa = _GEN_43[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_eff = _GEN_43[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_29_io_x_c = _GEN_43[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_ppn = _GEN_47[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_u = _GEN_47[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_ae = _GEN_47[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_sw = _GEN_47[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_sx = _GEN_47[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_sr = _GEN_47[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_pw = _GEN_47[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_px = _GEN_47[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_pr = _GEN_47[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_ppp = _GEN_47[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_pal = _GEN_47[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_paa = _GEN_47[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_eff = _GEN_47[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_30_io_x_c = _GEN_47[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_ppn = _GEN_51[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_u = _GEN_51[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_ae = _GEN_51[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_sw = _GEN_51[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_sx = _GEN_51[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_sr = _GEN_51[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_pw = _GEN_51[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_px = _GEN_51[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_pr = _GEN_51[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_ppp = _GEN_51[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_pal = _GEN_51[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_paa = _GEN_51[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_eff = _GEN_51[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_31_io_x_c = _GEN_51[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_ppn = _GEN_55[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_u = _GEN_55[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_ae = _GEN_55[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_sw = _GEN_55[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_sx = _GEN_55[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_sr = _GEN_55[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_pw = _GEN_55[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_px = _GEN_55[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_pr = _GEN_55[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_ppp = _GEN_55[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_pal = _GEN_55[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_paa = _GEN_55[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_eff = _GEN_55[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_32_io_x_c = _GEN_55[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_ppn = _GEN_59[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_u = _GEN_59[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_ae = _GEN_59[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_sw = _GEN_59[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_sx = _GEN_59[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_sr = _GEN_59[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_pw = _GEN_59[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_px = _GEN_59[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_pr = _GEN_59[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_ppp = _GEN_59[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_pal = _GEN_59[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_paa = _GEN_59[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_eff = _GEN_59[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_33_io_x_c = _GEN_59[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_ppn = _GEN_63[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_u = _GEN_63[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_ae = _GEN_63[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_sw = _GEN_63[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_sx = _GEN_63[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_sr = _GEN_63[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_pw = _GEN_63[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_px = _GEN_63[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_pr = _GEN_63[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_ppp = _GEN_63[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_pal = _GEN_63[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_paa = _GEN_63[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_eff = _GEN_63[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_34_io_x_c = _GEN_63[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_u = superpage_entries_0_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_ae = superpage_entries_0_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_sw = superpage_entries_0_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_sx = superpage_entries_0_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_sr = superpage_entries_0_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_pw = superpage_entries_0_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_px = superpage_entries_0_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_pr = superpage_entries_0_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_ppp = superpage_entries_0_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_35_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_u = superpage_entries_1_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_ae = superpage_entries_1_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_sw = superpage_entries_1_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_sx = superpage_entries_1_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_sr = superpage_entries_1_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_pw = superpage_entries_1_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_px = superpage_entries_1_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_pr = superpage_entries_1_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_ppp = superpage_entries_1_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_36_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_u = superpage_entries_2_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_ae = superpage_entries_2_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_sw = superpage_entries_2_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_sx = superpage_entries_2_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_sr = superpage_entries_2_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_pw = superpage_entries_2_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_px = superpage_entries_2_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_pr = superpage_entries_2_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_ppp = superpage_entries_2_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_37_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_u = superpage_entries_3_data_0[14]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_ae = superpage_entries_3_data_0[12]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_sw = superpage_entries_3_data_0[11]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_sx = superpage_entries_3_data_0[10]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_sr = superpage_entries_3_data_0[9]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_pw = superpage_entries_3_data_0[8]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_px = superpage_entries_3_data_0[7]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_pr = superpage_entries_3_data_0[6]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_ppp = superpage_entries_3_data_0[5]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 244:18]
  assign OptimizationBarrier_38_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 244:18]
  assign TLB_1_cov_read_addr = TLB_1_state;
  assign TLB_1_cov_read_data = TLB_1_cov[TLB_1_cov_read_addr]; // @[Coverage map for TLB_1]
  assign TLB_1_cov_write_data = 1'h1;
  assign TLB_1_cov_write_addr = TLB_1_state;
  assign TLB_1_cov_write_mask = 1'h1;
  assign TLB_1_cov_write_en = 1'h1;
  assign mux_cond_0 = sectored_entries_7_data_2[0];
  assign mux_cond_1 = ~sectored_entries_1_data_1[13];
  assign mux_cond_2 = ~sectored_entries_4_data_3[13];
  assign mux_cond_3 = ~sectored_entries_3_data_3[13];
  assign mux_cond_4 = sectored_entries_4_data_0[0];
  assign mux_cond_5 = sectored_entries_0_data_1[0];
  assign mux_cond_6 = sectored_entries_0_data_0[0];
  assign mux_cond_7 = sectored_entries_4_data_3[0];
  assign mux_cond_8 = sectored_entries_1_data_3[0];
  assign mux_cond_9 = sectored_entries_2_data_1[0];
  assign mux_cond_10 = ~sectored_entries_6_data_1[13];
  assign mux_cond_11 = ~sectored_entries_1_data_0[13];
  assign mux_cond_12 = sectored_entries_6_data_2[0];
  assign mux_cond_13 = ~sectored_entries_4_data_1[13];
  assign mux_cond_14 = sectored_entries_6_data_0[0];
  assign mux_cond_15 = sectored_entries_7_data_0[0];
  assign mux_cond_16 = sectored_entries_2_data_2[0];
  assign mux_cond_17 = sectored_entries_7_data_3[0];
  assign mux_cond_18 = ~sectored_entries_2_data_1[13];
  assign mux_cond_19 = sectored_entries_4_data_2[0];
  assign mux_cond_20 = ~sectored_entries_1_data_2[13];
  assign mux_cond_21 = ~superpage_entries_1_data_0[13];
  assign mux_cond_22 = ~sectored_entries_2_data_2[13];
  assign mux_cond_23 = ~sectored_entries_7_data_2[13];
  assign mux_cond_24 = ~sectored_entries_6_data_2[13];
  assign mux_cond_25 = ~sectored_entries_3_data_0[13];
  assign mux_cond_26 = sectored_entries_5_data_1[0];
  assign mux_cond_27 = sectored_entries_5_data_3[0];
  assign mux_cond_28 = ~sectored_entries_5_data_2[13];
  assign mux_cond_29 = sectored_entries_6_data_3[0];
  assign mux_cond_30 = ~sectored_entries_3_data_2[13];
  assign mux_cond_31 = ~sectored_entries_3_data_1[13];
  assign mux_cond_32 = sectored_entries_3_data_2[0];
  assign mux_cond_33 = ~sectored_entries_6_data_0[13];
  assign mux_cond_34 = sectored_entries_1_data_1[0];
  assign mux_cond_35 = ~sectored_entries_0_data_1[13];
  assign mux_cond_36 = sectored_entries_6_data_1[0];
  assign mux_cond_37 = sectored_entries_3_data_3[0];
  assign mux_cond_38 = ~sectored_entries_0_data_0[13];
  assign mux_cond_39 = sectored_entries_1_data_0[0];
  assign mux_cond_40 = ~sectored_entries_2_data_3[13];
  assign mux_cond_41 = sectored_entries_5_data_2[0];
  assign mux_cond_42 = sectored_entries_7_data_1[0];
  assign mux_cond_43 = ~sectored_entries_7_data_1[13];
  assign mux_cond_44 = sectored_entries_0_data_2[0];
  assign mux_cond_45 = sectored_entries_0_data_3[0];
  assign mux_cond_46 = ~sectored_entries_6_data_3[13];
  assign mux_cond_47 = sectored_entries_3_data_0[0];
  assign mux_cond_48 = ~sectored_entries_0_data_3[13];
  assign mux_cond_49 = sectored_entries_1_data_2[0];
  assign mux_cond_50 = sectored_entries_2_data_3[0];
  assign mux_cond_51 = sectored_entries_5_data_0[0];
  assign mux_cond_52 = ~sectored_entries_5_data_1[13];
  assign mux_cond_53 = ~sectored_entries_2_data_0[13];
  assign mux_cond_54 = ~sectored_entries_7_data_0[13];
  assign mux_cond_55 = ~sectored_entries_5_data_0[13];
  assign mux_cond_56 = ~sectored_entries_0_data_2[13];
  assign mux_cond_57 = ~superpage_entries_3_data_0[13];
  assign mux_cond_58 = ~special_entry_data_0[13];
  assign mux_cond_59 = sectored_entries_3_data_1[0];
  assign mux_cond_60 = sectored_entries_2_data_0[0];
  assign mux_cond_61 = ~sectored_entries_4_data_2[13];
  assign mux_cond_62 = ~sectored_entries_1_data_3[13];
  assign mux_cond_63 = ~superpage_entries_0_data_0[13];
  assign mux_cond_64 = sectored_entries_4_data_1[0];
  assign mux_cond_65 = ~sectored_entries_5_data_3[13];
  assign mux_cond_66 = ~superpage_entries_2_data_0[13];
  assign mux_cond_67 = ~sectored_entries_4_data_0[13];
  assign mux_cond_68 = ~sectored_entries_7_data_3[13];
  assign state_shl = {state, 2'h0};
  assign state_pad = {16'h0,state_shl};
  assign r_sectored_repl_addr_shl = r_sectored_repl_addr;
  assign r_sectored_repl_addr_pad = {17'h0,r_sectored_repl_addr_shl};
  assign r_superpage_repl_addr_shl = {r_superpage_repl_addr, 14'h0};
  assign r_superpage_repl_addr_pad = {4'h0,r_superpage_repl_addr_shl};
  assign r_sectored_hit_addr_shl = {r_sectored_hit_addr, 1'h0};
  assign r_sectored_hit_addr_pad = {16'h0,r_sectored_hit_addr_shl};
  assign special_entry_valid_0_shl = {special_entry_valid_0, 18'h0};
  assign special_entry_valid_0_pad = {1'h0,special_entry_valid_0_shl};
  assign r_sectored_hit_shl = {r_sectored_hit, 4'h0};
  assign r_sectored_hit_pad = {15'h0,r_sectored_hit_shl};
  assign special_entry_level_shl = {special_entry_level, 11'h0};
  assign special_entry_level_pad = {7'h0,special_entry_level_shl};
  assign mux_cond_0_shl = {mux_cond_0, 18'h0};
  assign mux_cond_0_pad = {1'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 8'h0};
  assign mux_cond_1_pad = {11'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 3'h0};
  assign mux_cond_2_pad = {16'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 18'h0};
  assign mux_cond_3_pad = {1'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 9'h0};
  assign mux_cond_4_pad = {10'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 12'h0};
  assign mux_cond_5_pad = {7'h0,mux_cond_5_shl};
  assign mux_cond_6_shl = {mux_cond_6, 12'h0};
  assign mux_cond_6_pad = {7'h0,mux_cond_6_shl};
  assign mux_cond_7_shl = {mux_cond_7, 6'h0};
  assign mux_cond_7_pad = {13'h0,mux_cond_7_shl};
  assign mux_cond_8_shl = {mux_cond_8, 1'h0};
  assign mux_cond_8_pad = {18'h0,mux_cond_8_shl};
  assign mux_cond_9_shl = {mux_cond_9, 17'h0};
  assign mux_cond_9_pad = {2'h0,mux_cond_9_shl};
  assign mux_cond_10_shl = {mux_cond_10, 5'h0};
  assign mux_cond_10_pad = {14'h0,mux_cond_10_shl};
  assign mux_cond_11_shl = mux_cond_11;
  assign mux_cond_11_pad = {19'h0,mux_cond_11_shl};
  assign mux_cond_12_shl = {mux_cond_12, 12'h0};
  assign mux_cond_12_pad = {7'h0,mux_cond_12_shl};
  assign mux_cond_13_shl = {mux_cond_13, 15'h0};
  assign mux_cond_13_pad = {4'h0,mux_cond_13_shl};
  assign mux_cond_14_shl = {mux_cond_14, 17'h0};
  assign mux_cond_14_pad = {2'h0,mux_cond_14_shl};
  assign mux_cond_15_shl = {mux_cond_15, 13'h0};
  assign mux_cond_15_pad = {6'h0,mux_cond_15_shl};
  assign mux_cond_16_shl = {mux_cond_16, 18'h0};
  assign mux_cond_16_pad = {1'h0,mux_cond_16_shl};
  assign mux_cond_17_shl = {mux_cond_17, 4'h0};
  assign mux_cond_17_pad = {15'h0,mux_cond_17_shl};
  assign mux_cond_18_shl = {mux_cond_18, 4'h0};
  assign mux_cond_18_pad = {15'h0,mux_cond_18_shl};
  assign mux_cond_19_shl = {mux_cond_19, 19'h0};
  assign mux_cond_19_pad = mux_cond_19_shl;
  assign mux_cond_20_shl = {mux_cond_20, 12'h0};
  assign mux_cond_20_pad = {7'h0,mux_cond_20_shl};
  assign mux_cond_21_shl = {mux_cond_21, 6'h0};
  assign mux_cond_21_pad = {13'h0,mux_cond_21_shl};
  assign mux_cond_22_shl = {mux_cond_22, 11'h0};
  assign mux_cond_22_pad = {8'h0,mux_cond_22_shl};
  assign mux_cond_23_shl = mux_cond_23;
  assign mux_cond_23_pad = {19'h0,mux_cond_23_shl};
  assign mux_cond_24_shl = mux_cond_24;
  assign mux_cond_24_pad = {19'h0,mux_cond_24_shl};
  assign mux_cond_25_shl = {mux_cond_25, 16'h0};
  assign mux_cond_25_pad = {3'h0,mux_cond_25_shl};
  assign mux_cond_26_shl = {mux_cond_26, 16'h0};
  assign mux_cond_26_pad = {3'h0,mux_cond_26_shl};
  assign mux_cond_27_shl = {mux_cond_27, 4'h0};
  assign mux_cond_27_pad = {15'h0,mux_cond_27_shl};
  assign mux_cond_28_shl = {mux_cond_28, 16'h0};
  assign mux_cond_28_pad = {3'h0,mux_cond_28_shl};
  assign mux_cond_29_shl = {mux_cond_29, 5'h0};
  assign mux_cond_29_pad = {14'h0,mux_cond_29_shl};
  assign mux_cond_30_shl = {mux_cond_30, 11'h0};
  assign mux_cond_30_pad = {8'h0,mux_cond_30_shl};
  assign mux_cond_31_shl = {mux_cond_31, 18'h0};
  assign mux_cond_31_pad = {1'h0,mux_cond_31_shl};
  assign mux_cond_32_shl = {mux_cond_32, 2'h0};
  assign mux_cond_32_pad = {17'h0,mux_cond_32_shl};
  assign mux_cond_33_shl = {mux_cond_33, 15'h0};
  assign mux_cond_33_pad = {4'h0,mux_cond_33_shl};
  assign mux_cond_34_shl = {mux_cond_34, 15'h0};
  assign mux_cond_34_pad = {4'h0,mux_cond_34_shl};
  assign mux_cond_35_shl = {mux_cond_35, 7'h0};
  assign mux_cond_35_pad = {12'h0,mux_cond_35_shl};
  assign mux_cond_36_shl = {mux_cond_36, 9'h0};
  assign mux_cond_36_pad = {10'h0,mux_cond_36_shl};
  assign mux_cond_37_shl = {mux_cond_37, 15'h0};
  assign mux_cond_37_pad = {4'h0,mux_cond_37_shl};
  assign mux_cond_38_shl = mux_cond_38;
  assign mux_cond_38_pad = {19'h0,mux_cond_38_shl};
  assign mux_cond_39_shl = {mux_cond_39, 12'h0};
  assign mux_cond_39_pad = {7'h0,mux_cond_39_shl};
  assign mux_cond_40_shl = {mux_cond_40, 15'h0};
  assign mux_cond_40_pad = {4'h0,mux_cond_40_shl};
  assign mux_cond_41_shl = {mux_cond_41, 13'h0};
  assign mux_cond_41_pad = {6'h0,mux_cond_41_shl};
  assign mux_cond_42_shl = {mux_cond_42, 7'h0};
  assign mux_cond_42_pad = {12'h0,mux_cond_42_shl};
  assign mux_cond_43_shl = {mux_cond_43, 2'h0};
  assign mux_cond_43_pad = {17'h0,mux_cond_43_shl};
  assign mux_cond_44_shl = {mux_cond_44, 6'h0};
  assign mux_cond_44_pad = {13'h0,mux_cond_44_shl};
  assign mux_cond_45_shl = {mux_cond_45, 8'h0};
  assign mux_cond_45_pad = {11'h0,mux_cond_45_shl};
  assign mux_cond_46_shl = {mux_cond_46, 13'h0};
  assign mux_cond_46_pad = {6'h0,mux_cond_46_shl};
  assign mux_cond_47_shl = {mux_cond_47, 19'h0};
  assign mux_cond_47_pad = mux_cond_47_shl;
  assign mux_cond_48_shl = {mux_cond_48, 10'h0};
  assign mux_cond_48_pad = {9'h0,mux_cond_48_shl};
  assign mux_cond_49_shl = {mux_cond_49, 2'h0};
  assign mux_cond_49_pad = {17'h0,mux_cond_49_shl};
  assign mux_cond_50_shl = {mux_cond_50, 6'h0};
  assign mux_cond_50_pad = {13'h0,mux_cond_50_shl};
  assign mux_cond_51_shl = {mux_cond_51, 2'h0};
  assign mux_cond_51_pad = {17'h0,mux_cond_51_shl};
  assign mux_cond_52_shl = {mux_cond_52, 8'h0};
  assign mux_cond_52_pad = {11'h0,mux_cond_52_shl};
  assign mux_cond_53_shl = {mux_cond_53, 11'h0};
  assign mux_cond_53_pad = {8'h0,mux_cond_53_shl};
  assign mux_cond_54_shl = {mux_cond_54, 8'h0};
  assign mux_cond_54_pad = {11'h0,mux_cond_54_shl};
  assign mux_cond_55_shl = {mux_cond_55, 12'h0};
  assign mux_cond_55_pad = {7'h0,mux_cond_55_shl};
  assign mux_cond_56_shl = {mux_cond_56, 10'h0};
  assign mux_cond_56_pad = {9'h0,mux_cond_56_shl};
  assign mux_cond_57_shl = {mux_cond_57, 3'h0};
  assign mux_cond_57_pad = {16'h0,mux_cond_57_shl};
  assign mux_cond_58_shl = mux_cond_58;
  assign mux_cond_58_pad = {19'h0,mux_cond_58_shl};
  assign mux_cond_59_shl = {mux_cond_59, 11'h0};
  assign mux_cond_59_pad = {8'h0,mux_cond_59_shl};
  assign mux_cond_60_shl = {mux_cond_60, 3'h0};
  assign mux_cond_60_pad = {16'h0,mux_cond_60_shl};
  assign mux_cond_61_shl = {mux_cond_61, 13'h0};
  assign mux_cond_61_pad = {6'h0,mux_cond_61_shl};
  assign mux_cond_62_shl = {mux_cond_62, 8'h0};
  assign mux_cond_62_pad = {11'h0,mux_cond_62_shl};
  assign mux_cond_63_shl = mux_cond_63;
  assign mux_cond_63_pad = {19'h0,mux_cond_63_shl};
  assign mux_cond_64_shl = {mux_cond_64, 6'h0};
  assign mux_cond_64_pad = {13'h0,mux_cond_64_shl};
  assign mux_cond_65_shl = {mux_cond_65, 13'h0};
  assign mux_cond_65_pad = {6'h0,mux_cond_65_shl};
  assign mux_cond_66_shl = {mux_cond_66, 4'h0};
  assign mux_cond_66_pad = {15'h0,mux_cond_66_shl};
  assign mux_cond_67_shl = {mux_cond_67, 10'h0};
  assign mux_cond_67_pad = {9'h0,mux_cond_67_shl};
  assign mux_cond_68_shl = {mux_cond_68, 15'h0};
  assign mux_cond_68_pad = {4'h0,mux_cond_68_shl};
  assign superpage_entries_2_level_shl = {superpage_entries_2_level, 16'h0};
  assign superpage_entries_2_level_pad = {2'h0,superpage_entries_2_level_shl};
  assign sectored_entries_7_valid_3_shl = {sectored_entries_7_valid_3, 14'h0};
  assign sectored_entries_7_valid_3_pad = {5'h0,sectored_entries_7_valid_3_shl};
  assign superpage_entries_1_level_shl = {superpage_entries_1_level, 16'h0};
  assign superpage_entries_1_level_pad = {2'h0,superpage_entries_1_level_shl};
  assign superpage_entries_1_valid_0_shl = {superpage_entries_1_valid_0, 11'h0};
  assign superpage_entries_1_valid_0_pad = {8'h0,superpage_entries_1_valid_0_shl};
  assign sectored_entries_3_valid_0_shl = {sectored_entries_3_valid_0, 18'h0};
  assign sectored_entries_3_valid_0_pad = {1'h0,sectored_entries_3_valid_0_shl};
  assign sectored_entries_1_valid_3_shl = {sectored_entries_1_valid_3, 14'h0};
  assign sectored_entries_1_valid_3_pad = {5'h0,sectored_entries_1_valid_3_shl};
  assign sectored_entries_6_valid_3_shl = {sectored_entries_6_valid_3, 14'h0};
  assign sectored_entries_6_valid_3_pad = {5'h0,sectored_entries_6_valid_3_shl};
  assign sectored_entries_1_valid_0_shl = {sectored_entries_1_valid_0, 18'h0};
  assign sectored_entries_1_valid_0_pad = {1'h0,sectored_entries_1_valid_0_shl};
  assign sectored_entries_2_valid_0_shl = {sectored_entries_2_valid_0, 18'h0};
  assign sectored_entries_2_valid_0_pad = {1'h0,sectored_entries_2_valid_0_shl};
  assign sectored_entries_3_valid_1_shl = {sectored_entries_3_valid_1, 14'h0};
  assign sectored_entries_3_valid_1_pad = {5'h0,sectored_entries_3_valid_1_shl};
  assign sectored_entries_5_valid_3_shl = {sectored_entries_5_valid_3, 14'h0};
  assign sectored_entries_5_valid_3_pad = {5'h0,sectored_entries_5_valid_3_shl};
  assign superpage_entries_3_valid_0_shl = {superpage_entries_3_valid_0, 11'h0};
  assign superpage_entries_3_valid_0_pad = {8'h0,superpage_entries_3_valid_0_shl};
  assign sectored_entries_5_valid_1_shl = {sectored_entries_5_valid_1, 14'h0};
  assign sectored_entries_5_valid_1_pad = {5'h0,sectored_entries_5_valid_1_shl};
  assign sectored_entries_0_valid_3_shl = {sectored_entries_0_valid_3, 14'h0};
  assign sectored_entries_0_valid_3_pad = {5'h0,sectored_entries_0_valid_3_shl};
  assign sectored_entries_6_valid_0_shl = {sectored_entries_6_valid_0, 18'h0};
  assign sectored_entries_6_valid_0_pad = {1'h0,sectored_entries_6_valid_0_shl};
  assign sectored_entries_0_valid_0_shl = {sectored_entries_0_valid_0, 18'h0};
  assign sectored_entries_0_valid_0_pad = {1'h0,sectored_entries_0_valid_0_shl};
  assign sectored_entries_4_valid_2_shl = {sectored_entries_4_valid_2, 16'h0};
  assign sectored_entries_4_valid_2_pad = {3'h0,sectored_entries_4_valid_2_shl};
  assign superpage_entries_2_valid_0_shl = {superpage_entries_2_valid_0, 11'h0};
  assign superpage_entries_2_valid_0_pad = {8'h0,superpage_entries_2_valid_0_shl};
  assign sectored_entries_2_valid_1_shl = {sectored_entries_2_valid_1, 14'h0};
  assign sectored_entries_2_valid_1_pad = {5'h0,sectored_entries_2_valid_1_shl};
  assign superpage_entries_0_level_shl = {superpage_entries_0_level, 16'h0};
  assign superpage_entries_0_level_pad = {2'h0,superpage_entries_0_level_shl};
  assign sectored_entries_1_valid_1_shl = {sectored_entries_1_valid_1, 14'h0};
  assign sectored_entries_1_valid_1_pad = {5'h0,sectored_entries_1_valid_1_shl};
  assign sectored_entries_4_valid_3_shl = {sectored_entries_4_valid_3, 14'h0};
  assign sectored_entries_4_valid_3_pad = {5'h0,sectored_entries_4_valid_3_shl};
  assign sectored_entries_0_valid_1_shl = {sectored_entries_0_valid_1, 14'h0};
  assign sectored_entries_0_valid_1_pad = {5'h0,sectored_entries_0_valid_1_shl};
  assign sectored_entries_4_valid_0_shl = {sectored_entries_4_valid_0, 18'h0};
  assign sectored_entries_4_valid_0_pad = {1'h0,sectored_entries_4_valid_0_shl};
  assign sectored_entries_0_valid_2_shl = {sectored_entries_0_valid_2, 16'h0};
  assign sectored_entries_0_valid_2_pad = {3'h0,sectored_entries_0_valid_2_shl};
  assign sectored_entries_1_valid_2_shl = {sectored_entries_1_valid_2, 16'h0};
  assign sectored_entries_1_valid_2_pad = {3'h0,sectored_entries_1_valid_2_shl};
  assign sectored_entries_2_valid_2_shl = {sectored_entries_2_valid_2, 16'h0};
  assign sectored_entries_2_valid_2_pad = {3'h0,sectored_entries_2_valid_2_shl};
  assign sectored_entries_7_valid_0_shl = {sectored_entries_7_valid_0, 18'h0};
  assign sectored_entries_7_valid_0_pad = {1'h0,sectored_entries_7_valid_0_shl};
  assign sectored_entries_5_valid_2_shl = {sectored_entries_5_valid_2, 16'h0};
  assign sectored_entries_5_valid_2_pad = {3'h0,sectored_entries_5_valid_2_shl};
  assign sectored_entries_7_valid_2_shl = {sectored_entries_7_valid_2, 16'h0};
  assign sectored_entries_7_valid_2_pad = {3'h0,sectored_entries_7_valid_2_shl};
  assign sectored_entries_4_valid_1_shl = {sectored_entries_4_valid_1, 14'h0};
  assign sectored_entries_4_valid_1_pad = {5'h0,sectored_entries_4_valid_1_shl};
  assign sectored_entries_5_valid_0_shl = {sectored_entries_5_valid_0, 18'h0};
  assign sectored_entries_5_valid_0_pad = {1'h0,sectored_entries_5_valid_0_shl};
  assign sectored_entries_7_valid_1_shl = {sectored_entries_7_valid_1, 14'h0};
  assign sectored_entries_7_valid_1_pad = {5'h0,sectored_entries_7_valid_1_shl};
  assign superpage_entries_3_level_shl = {superpage_entries_3_level, 16'h0};
  assign superpage_entries_3_level_pad = {2'h0,superpage_entries_3_level_shl};
  assign sectored_entries_3_valid_3_shl = {sectored_entries_3_valid_3, 14'h0};
  assign sectored_entries_3_valid_3_pad = {5'h0,sectored_entries_3_valid_3_shl};
  assign sectored_entries_2_valid_3_shl = {sectored_entries_2_valid_3, 14'h0};
  assign sectored_entries_2_valid_3_pad = {5'h0,sectored_entries_2_valid_3_shl};
  assign superpage_entries_0_valid_0_shl = {superpage_entries_0_valid_0, 11'h0};
  assign superpage_entries_0_valid_0_pad = {8'h0,superpage_entries_0_valid_0_shl};
  assign sectored_entries_6_valid_1_shl = {sectored_entries_6_valid_1, 14'h0};
  assign sectored_entries_6_valid_1_pad = {5'h0,sectored_entries_6_valid_1_shl};
  assign sectored_entries_3_valid_2_shl = {sectored_entries_3_valid_2, 16'h0};
  assign sectored_entries_3_valid_2_pad = {3'h0,sectored_entries_3_valid_2_shl};
  assign sectored_entries_6_valid_2_shl = {sectored_entries_6_valid_2, 16'h0};
  assign sectored_entries_6_valid_2_pad = {3'h0,sectored_entries_6_valid_2_shl};
  assign TLB_1_xor64 = r_sectored_repl_addr_pad ^ r_superpage_repl_addr_pad;
  assign TLB_1_xor31 = state_pad ^ TLB_1_xor64;
  assign TLB_1_xor65 = r_sectored_hit_addr_pad ^ special_entry_valid_0_pad;
  assign TLB_1_xor66 = r_sectored_hit_pad ^ special_entry_level_pad;
  assign TLB_1_xor32 = TLB_1_xor65 ^ TLB_1_xor66;
  assign TLB_1_xor15 = TLB_1_xor31 ^ TLB_1_xor32;
  assign TLB_1_xor68 = mux_cond_1_pad ^ mux_cond_2_pad;
  assign TLB_1_xor33 = mux_cond_0_pad ^ TLB_1_xor68;
  assign TLB_1_xor69 = mux_cond_3_pad ^ mux_cond_4_pad;
  assign TLB_1_xor70 = mux_cond_5_pad ^ mux_cond_6_pad;
  assign TLB_1_xor34 = TLB_1_xor69 ^ TLB_1_xor70;
  assign TLB_1_xor16 = TLB_1_xor33 ^ TLB_1_xor34;
  assign TLB_1_xor7 = TLB_1_xor15 ^ TLB_1_xor16;
  assign TLB_1_xor72 = mux_cond_8_pad ^ mux_cond_9_pad;
  assign TLB_1_xor35 = mux_cond_7_pad ^ TLB_1_xor72;
  assign TLB_1_xor73 = mux_cond_10_pad ^ mux_cond_11_pad;
  assign TLB_1_xor74 = mux_cond_12_pad ^ mux_cond_13_pad;
  assign TLB_1_xor36 = TLB_1_xor73 ^ TLB_1_xor74;
  assign TLB_1_xor17 = TLB_1_xor35 ^ TLB_1_xor36;
  assign TLB_1_xor75 = mux_cond_14_pad ^ mux_cond_15_pad;
  assign TLB_1_xor76 = mux_cond_16_pad ^ mux_cond_17_pad;
  assign TLB_1_xor37 = TLB_1_xor75 ^ TLB_1_xor76;
  assign TLB_1_xor77 = mux_cond_18_pad ^ mux_cond_19_pad;
  assign TLB_1_xor78 = mux_cond_20_pad ^ mux_cond_21_pad;
  assign TLB_1_xor38 = TLB_1_xor77 ^ TLB_1_xor78;
  assign TLB_1_xor18 = TLB_1_xor37 ^ TLB_1_xor38;
  assign TLB_1_xor8 = TLB_1_xor17 ^ TLB_1_xor18;
  assign TLB_1_xor3 = TLB_1_xor7 ^ TLB_1_xor8;
  assign TLB_1_xor80 = mux_cond_23_pad ^ mux_cond_24_pad;
  assign TLB_1_xor39 = mux_cond_22_pad ^ TLB_1_xor80;
  assign TLB_1_xor81 = mux_cond_25_pad ^ mux_cond_26_pad;
  assign TLB_1_xor82 = mux_cond_27_pad ^ mux_cond_28_pad;
  assign TLB_1_xor40 = TLB_1_xor81 ^ TLB_1_xor82;
  assign TLB_1_xor19 = TLB_1_xor39 ^ TLB_1_xor40;
  assign TLB_1_xor84 = mux_cond_30_pad ^ mux_cond_31_pad;
  assign TLB_1_xor41 = mux_cond_29_pad ^ TLB_1_xor84;
  assign TLB_1_xor85 = mux_cond_32_pad ^ mux_cond_33_pad;
  assign TLB_1_xor86 = mux_cond_34_pad ^ mux_cond_35_pad;
  assign TLB_1_xor42 = TLB_1_xor85 ^ TLB_1_xor86;
  assign TLB_1_xor20 = TLB_1_xor41 ^ TLB_1_xor42;
  assign TLB_1_xor9 = TLB_1_xor19 ^ TLB_1_xor20;
  assign TLB_1_xor88 = mux_cond_37_pad ^ mux_cond_38_pad;
  assign TLB_1_xor43 = mux_cond_36_pad ^ TLB_1_xor88;
  assign TLB_1_xor89 = mux_cond_39_pad ^ mux_cond_40_pad;
  assign TLB_1_xor90 = mux_cond_41_pad ^ mux_cond_42_pad;
  assign TLB_1_xor44 = TLB_1_xor89 ^ TLB_1_xor90;
  assign TLB_1_xor21 = TLB_1_xor43 ^ TLB_1_xor44;
  assign TLB_1_xor91 = mux_cond_43_pad ^ mux_cond_44_pad;
  assign TLB_1_xor92 = mux_cond_45_pad ^ mux_cond_46_pad;
  assign TLB_1_xor45 = TLB_1_xor91 ^ TLB_1_xor92;
  assign TLB_1_xor93 = mux_cond_47_pad ^ mux_cond_48_pad;
  assign TLB_1_xor94 = mux_cond_49_pad ^ mux_cond_50_pad;
  assign TLB_1_xor46 = TLB_1_xor93 ^ TLB_1_xor94;
  assign TLB_1_xor22 = TLB_1_xor45 ^ TLB_1_xor46;
  assign TLB_1_xor10 = TLB_1_xor21 ^ TLB_1_xor22;
  assign TLB_1_xor4 = TLB_1_xor9 ^ TLB_1_xor10;
  assign TLB_1_xor1 = TLB_1_xor3 ^ TLB_1_xor4;
  assign TLB_1_xor96 = mux_cond_52_pad ^ mux_cond_53_pad;
  assign TLB_1_xor47 = mux_cond_51_pad ^ TLB_1_xor96;
  assign TLB_1_xor97 = mux_cond_54_pad ^ mux_cond_55_pad;
  assign TLB_1_xor98 = mux_cond_56_pad ^ mux_cond_57_pad;
  assign TLB_1_xor48 = TLB_1_xor97 ^ TLB_1_xor98;
  assign TLB_1_xor23 = TLB_1_xor47 ^ TLB_1_xor48;
  assign TLB_1_xor100 = mux_cond_59_pad ^ mux_cond_60_pad;
  assign TLB_1_xor49 = mux_cond_58_pad ^ TLB_1_xor100;
  assign TLB_1_xor101 = mux_cond_61_pad ^ mux_cond_62_pad;
  assign TLB_1_xor102 = mux_cond_63_pad ^ mux_cond_64_pad;
  assign TLB_1_xor50 = TLB_1_xor101 ^ TLB_1_xor102;
  assign TLB_1_xor24 = TLB_1_xor49 ^ TLB_1_xor50;
  assign TLB_1_xor11 = TLB_1_xor23 ^ TLB_1_xor24;
  assign TLB_1_xor104 = mux_cond_66_pad ^ mux_cond_67_pad;
  assign TLB_1_xor51 = mux_cond_65_pad ^ TLB_1_xor104;
  assign TLB_1_xor105 = mux_cond_68_pad ^ superpage_entries_2_level_pad;
  assign TLB_1_xor106 = sectored_entries_7_valid_3_pad ^ superpage_entries_1_level_pad;
  assign TLB_1_xor52 = TLB_1_xor105 ^ TLB_1_xor106;
  assign TLB_1_xor25 = TLB_1_xor51 ^ TLB_1_xor52;
  assign TLB_1_xor107 = superpage_entries_1_valid_0_pad ^ sectored_entries_3_valid_0_pad;
  assign TLB_1_xor108 = sectored_entries_1_valid_3_pad ^ sectored_entries_6_valid_3_pad;
  assign TLB_1_xor53 = TLB_1_xor107 ^ TLB_1_xor108;
  assign TLB_1_xor109 = sectored_entries_1_valid_0_pad ^ sectored_entries_2_valid_0_pad;
  assign TLB_1_xor110 = sectored_entries_3_valid_1_pad ^ sectored_entries_5_valid_3_pad;
  assign TLB_1_xor54 = TLB_1_xor109 ^ TLB_1_xor110;
  assign TLB_1_xor26 = TLB_1_xor53 ^ TLB_1_xor54;
  assign TLB_1_xor12 = TLB_1_xor25 ^ TLB_1_xor26;
  assign TLB_1_xor5 = TLB_1_xor11 ^ TLB_1_xor12;
  assign TLB_1_xor112 = sectored_entries_5_valid_1_pad ^ sectored_entries_0_valid_3_pad;
  assign TLB_1_xor55 = superpage_entries_3_valid_0_pad ^ TLB_1_xor112;
  assign TLB_1_xor113 = sectored_entries_6_valid_0_pad ^ sectored_entries_0_valid_0_pad;
  assign TLB_1_xor114 = sectored_entries_4_valid_2_pad ^ superpage_entries_2_valid_0_pad;
  assign TLB_1_xor56 = TLB_1_xor113 ^ TLB_1_xor114;
  assign TLB_1_xor27 = TLB_1_xor55 ^ TLB_1_xor56;
  assign TLB_1_xor116 = superpage_entries_0_level_pad ^ sectored_entries_1_valid_1_pad;
  assign TLB_1_xor57 = sectored_entries_2_valid_1_pad ^ TLB_1_xor116;
  assign TLB_1_xor117 = sectored_entries_4_valid_3_pad ^ sectored_entries_0_valid_1_pad;
  assign TLB_1_xor118 = sectored_entries_4_valid_0_pad ^ sectored_entries_0_valid_2_pad;
  assign TLB_1_xor58 = TLB_1_xor117 ^ TLB_1_xor118;
  assign TLB_1_xor28 = TLB_1_xor57 ^ TLB_1_xor58;
  assign TLB_1_xor13 = TLB_1_xor27 ^ TLB_1_xor28;
  assign TLB_1_xor120 = sectored_entries_2_valid_2_pad ^ sectored_entries_7_valid_0_pad;
  assign TLB_1_xor59 = sectored_entries_1_valid_2_pad ^ TLB_1_xor120;
  assign TLB_1_xor121 = sectored_entries_5_valid_2_pad ^ sectored_entries_7_valid_2_pad;
  assign TLB_1_xor122 = sectored_entries_4_valid_1_pad ^ sectored_entries_5_valid_0_pad;
  assign TLB_1_xor60 = TLB_1_xor121 ^ TLB_1_xor122;
  assign TLB_1_xor29 = TLB_1_xor59 ^ TLB_1_xor60;
  assign TLB_1_xor123 = sectored_entries_7_valid_1_pad ^ superpage_entries_3_level_pad;
  assign TLB_1_xor124 = sectored_entries_3_valid_3_pad ^ sectored_entries_2_valid_3_pad;
  assign TLB_1_xor61 = TLB_1_xor123 ^ TLB_1_xor124;
  assign TLB_1_xor125 = superpage_entries_0_valid_0_pad ^ sectored_entries_6_valid_1_pad;
  assign TLB_1_xor126 = sectored_entries_3_valid_2_pad ^ sectored_entries_6_valid_2_pad;
  assign TLB_1_xor62 = TLB_1_xor125 ^ TLB_1_xor126;
  assign TLB_1_xor30 = TLB_1_xor61 ^ TLB_1_xor62;
  assign TLB_1_xor14 = TLB_1_xor29 ^ TLB_1_xor30;
  assign TLB_1_xor6 = TLB_1_xor13 ^ TLB_1_xor14;
  assign TLB_1_xor2 = TLB_1_xor5 ^ TLB_1_xor6;
  assign TLB_1_xor0 = TLB_1_xor1 ^ TLB_1_xor2;
  assign OptimizationBarrier_20_sum = TLB_1_covSum + OptimizationBarrier_20_io_covSum;
  assign OptimizationBarrier_21_sum = OptimizationBarrier_20_sum + OptimizationBarrier_21_io_covSum;
  assign OptimizationBarrier_35_sum = OptimizationBarrier_21_sum + OptimizationBarrier_35_io_covSum;
  assign OptimizationBarrier_6_sum = OptimizationBarrier_35_sum + OptimizationBarrier_6_io_covSum;
  assign OptimizationBarrier_16_sum = OptimizationBarrier_6_sum + OptimizationBarrier_16_io_covSum;
  assign OptimizationBarrier_12_sum = OptimizationBarrier_16_sum + OptimizationBarrier_12_io_covSum;
  assign OptimizationBarrier_9_sum = OptimizationBarrier_12_sum + OptimizationBarrier_9_io_covSum;
  assign OptimizationBarrier_8_sum = OptimizationBarrier_9_sum + OptimizationBarrier_8_io_covSum;
  assign OptimizationBarrier_2_sum = OptimizationBarrier_8_sum + OptimizationBarrier_2_io_covSum;
  assign OptimizationBarrier_25_sum = OptimizationBarrier_2_sum + OptimizationBarrier_25_io_covSum;
  assign OptimizationBarrier_23_sum = OptimizationBarrier_25_sum + OptimizationBarrier_23_io_covSum;
  assign OptimizationBarrier_27_sum = OptimizationBarrier_23_sum + OptimizationBarrier_27_io_covSum;
  assign OptimizationBarrier_30_sum = OptimizationBarrier_27_sum + OptimizationBarrier_30_io_covSum;
  assign OptimizationBarrier_1_sum = OptimizationBarrier_30_sum + OptimizationBarrier_1_io_covSum;
  assign OptimizationBarrier_18_sum = OptimizationBarrier_1_sum + OptimizationBarrier_18_io_covSum;
  assign OptimizationBarrier_31_sum = OptimizationBarrier_18_sum + OptimizationBarrier_31_io_covSum;
  assign OptimizationBarrier_19_sum = OptimizationBarrier_31_sum + OptimizationBarrier_19_io_covSum;
  assign OptimizationBarrier_37_sum = OptimizationBarrier_19_sum + OptimizationBarrier_37_io_covSum;
  assign OptimizationBarrier_28_sum = OptimizationBarrier_37_sum + OptimizationBarrier_28_io_covSum;
  assign OptimizationBarrier_33_sum = OptimizationBarrier_28_sum + OptimizationBarrier_33_io_covSum;
  assign OptimizationBarrier_4_sum = OptimizationBarrier_33_sum + OptimizationBarrier_4_io_covSum;
  assign OptimizationBarrier_38_sum = OptimizationBarrier_4_sum + OptimizationBarrier_38_io_covSum;
  assign pmp_sum = OptimizationBarrier_38_sum + pmp_io_covSum;
  assign OptimizationBarrier_sum = pmp_sum + OptimizationBarrier_io_covSum;
  assign OptimizationBarrier_34_sum = OptimizationBarrier_sum + OptimizationBarrier_34_io_covSum;
  assign OptimizationBarrier_24_sum = OptimizationBarrier_34_sum + OptimizationBarrier_24_io_covSum;
  assign OptimizationBarrier_22_sum = OptimizationBarrier_24_sum + OptimizationBarrier_22_io_covSum;
  assign OptimizationBarrier_10_sum = OptimizationBarrier_22_sum + OptimizationBarrier_10_io_covSum;
  assign OptimizationBarrier_3_sum = OptimizationBarrier_10_sum + OptimizationBarrier_3_io_covSum;
  assign OptimizationBarrier_5_sum = OptimizationBarrier_3_sum + OptimizationBarrier_5_io_covSum;
  assign OptimizationBarrier_36_sum = OptimizationBarrier_5_sum + OptimizationBarrier_36_io_covSum;
  assign OptimizationBarrier_17_sum = OptimizationBarrier_36_sum + OptimizationBarrier_17_io_covSum;
  assign OptimizationBarrier_15_sum = OptimizationBarrier_17_sum + OptimizationBarrier_15_io_covSum;
  assign OptimizationBarrier_29_sum = OptimizationBarrier_15_sum + OptimizationBarrier_29_io_covSum;
  assign OptimizationBarrier_32_sum = OptimizationBarrier_29_sum + OptimizationBarrier_32_io_covSum;
  assign OptimizationBarrier_7_sum = OptimizationBarrier_32_sum + OptimizationBarrier_7_io_covSum;
  assign OptimizationBarrier_14_sum = OptimizationBarrier_7_sum + OptimizationBarrier_14_io_covSum;
  assign OptimizationBarrier_26_sum = OptimizationBarrier_14_sum + OptimizationBarrier_26_io_covSum;
  assign OptimizationBarrier_11_sum = OptimizationBarrier_26_sum + OptimizationBarrier_11_io_covSum;
  assign OptimizationBarrier_13_sum = OptimizationBarrier_11_sum + OptimizationBarrier_13_io_covSum;
  assign io_covSum = OptimizationBarrier_13_sum;
  assign stopEn0 = io_sfence_valid & ~_T_2454;
  assign OptimizationBarrier_38_metaAssert_wire = OptimizationBarrier_38_metaAssert;
  assign OptimizationBarrier_2_metaAssert_wire = OptimizationBarrier_2_metaAssert;
  assign OptimizationBarrier_26_metaAssert_wire = OptimizationBarrier_26_metaAssert;
  assign OptimizationBarrier_metaAssert_wire = OptimizationBarrier_metaAssert;
  assign OptimizationBarrier_7_metaAssert_wire = OptimizationBarrier_7_metaAssert;
  assign OptimizationBarrier_37_metaAssert_wire = OptimizationBarrier_37_metaAssert;
  assign OptimizationBarrier_24_metaAssert_wire = OptimizationBarrier_24_metaAssert;
  assign OptimizationBarrier_17_metaAssert_wire = OptimizationBarrier_17_metaAssert;
  assign OptimizationBarrier_34_metaAssert_wire = OptimizationBarrier_34_metaAssert;
  assign OptimizationBarrier_21_metaAssert_wire = OptimizationBarrier_21_metaAssert;
  assign OptimizationBarrier_28_metaAssert_wire = OptimizationBarrier_28_metaAssert;
  assign OptimizationBarrier_16_metaAssert_wire = OptimizationBarrier_16_metaAssert;
  assign OptimizationBarrier_5_metaAssert_wire = OptimizationBarrier_5_metaAssert;
  assign OptimizationBarrier_8_metaAssert_wire = OptimizationBarrier_8_metaAssert;
  assign OptimizationBarrier_1_metaAssert_wire = OptimizationBarrier_1_metaAssert;
  assign OptimizationBarrier_4_metaAssert_wire = OptimizationBarrier_4_metaAssert;
  assign OptimizationBarrier_33_metaAssert_wire = OptimizationBarrier_33_metaAssert;
  assign OptimizationBarrier_30_metaAssert_wire = OptimizationBarrier_30_metaAssert;
  assign OptimizationBarrier_19_metaAssert_wire = OptimizationBarrier_19_metaAssert;
  assign OptimizationBarrier_20_metaAssert_wire = OptimizationBarrier_20_metaAssert;
  assign OptimizationBarrier_9_metaAssert_wire = OptimizationBarrier_9_metaAssert;
  assign OptimizationBarrier_29_metaAssert_wire = OptimizationBarrier_29_metaAssert;
  assign OptimizationBarrier_36_metaAssert_wire = OptimizationBarrier_36_metaAssert;
  assign OptimizationBarrier_31_metaAssert_wire = OptimizationBarrier_31_metaAssert;
  assign OptimizationBarrier_18_metaAssert_wire = OptimizationBarrier_18_metaAssert;
  assign OptimizationBarrier_12_metaAssert_wire = OptimizationBarrier_12_metaAssert;
  assign OptimizationBarrier_23_metaAssert_wire = OptimizationBarrier_23_metaAssert;
  assign OptimizationBarrier_32_metaAssert_wire = OptimizationBarrier_32_metaAssert;
  assign OptimizationBarrier_25_metaAssert_wire = OptimizationBarrier_25_metaAssert;
  assign OptimizationBarrier_6_metaAssert_wire = OptimizationBarrier_6_metaAssert;
  assign pmp_metaAssert_wire = pmp_metaAssert;
  assign OptimizationBarrier_27_metaAssert_wire = OptimizationBarrier_27_metaAssert;
  assign OptimizationBarrier_3_metaAssert_wire = OptimizationBarrier_3_metaAssert;
  assign OptimizationBarrier_14_metaAssert_wire = OptimizationBarrier_14_metaAssert;
  assign OptimizationBarrier_11_metaAssert_wire = OptimizationBarrier_11_metaAssert;
  assign OptimizationBarrier_15_metaAssert_wire = OptimizationBarrier_15_metaAssert;
  assign OptimizationBarrier_13_metaAssert_wire = OptimizationBarrier_13_metaAssert;
  assign OptimizationBarrier_22_metaAssert_wire = OptimizationBarrier_22_metaAssert;
  assign OptimizationBarrier_35_metaAssert_wire = OptimizationBarrier_35_metaAssert;
  assign OptimizationBarrier_10_metaAssert_wire = OptimizationBarrier_10_metaAssert;
  assign TLB_1_or15 = stopEn0 | OptimizationBarrier_33_metaAssert_wire;
  assign TLB_1_or34 = OptimizationBarrier_5_metaAssert_wire | OptimizationBarrier_20_metaAssert_wire;
  assign TLB_1_or16 = OptimizationBarrier_7_metaAssert_wire | TLB_1_or34;
  assign TLB_1_or7 = TLB_1_or15 | TLB_1_or16;
  assign TLB_1_or17 = OptimizationBarrier_22_metaAssert_wire | OptimizationBarrier_14_metaAssert_wire;
  assign TLB_1_or38 = OptimizationBarrier_metaAssert_wire | OptimizationBarrier_31_metaAssert_wire;
  assign TLB_1_or18 = OptimizationBarrier_2_metaAssert_wire | TLB_1_or38;
  assign TLB_1_or8 = TLB_1_or17 | TLB_1_or18;
  assign TLB_1_or3 = TLB_1_or7 | TLB_1_or8;
  assign TLB_1_or19 = OptimizationBarrier_18_metaAssert_wire | OptimizationBarrier_24_metaAssert_wire;
  assign TLB_1_or42 = OptimizationBarrier_25_metaAssert_wire | OptimizationBarrier_13_metaAssert_wire;
  assign TLB_1_or20 = OptimizationBarrier_10_metaAssert_wire | TLB_1_or42;
  assign TLB_1_or9 = TLB_1_or19 | TLB_1_or20;
  assign TLB_1_or21 = OptimizationBarrier_36_metaAssert_wire | OptimizationBarrier_34_metaAssert_wire;
  assign TLB_1_or46 = OptimizationBarrier_8_metaAssert_wire | OptimizationBarrier_21_metaAssert_wire;
  assign TLB_1_or22 = OptimizationBarrier_16_metaAssert_wire | TLB_1_or46;
  assign TLB_1_or10 = TLB_1_or21 | TLB_1_or22;
  assign TLB_1_or4 = TLB_1_or9 | TLB_1_or10;
  assign TLB_1_or1 = TLB_1_or3 | TLB_1_or4;
  assign TLB_1_or23 = OptimizationBarrier_12_metaAssert_wire | OptimizationBarrier_30_metaAssert_wire;
  assign TLB_1_or50 = OptimizationBarrier_27_metaAssert_wire | OptimizationBarrier_32_metaAssert_wire;
  assign TLB_1_or24 = pmp_metaAssert_wire | TLB_1_or50;
  assign TLB_1_or11 = TLB_1_or23 | TLB_1_or24;
  assign TLB_1_or25 = OptimizationBarrier_29_metaAssert_wire | OptimizationBarrier_1_metaAssert_wire;
  assign TLB_1_or54 = OptimizationBarrier_3_metaAssert_wire | OptimizationBarrier_38_metaAssert_wire;
  assign TLB_1_or26 = OptimizationBarrier_9_metaAssert_wire | TLB_1_or54;
  assign TLB_1_or12 = TLB_1_or25 | TLB_1_or26;
  assign TLB_1_or5 = TLB_1_or11 | TLB_1_or12;
  assign TLB_1_or27 = OptimizationBarrier_4_metaAssert_wire | OptimizationBarrier_6_metaAssert_wire;
  assign TLB_1_or58 = OptimizationBarrier_26_metaAssert_wire | OptimizationBarrier_19_metaAssert_wire;
  assign TLB_1_or28 = OptimizationBarrier_37_metaAssert_wire | TLB_1_or58;
  assign TLB_1_or13 = TLB_1_or27 | TLB_1_or28;
  assign TLB_1_or60 = OptimizationBarrier_11_metaAssert_wire | OptimizationBarrier_15_metaAssert_wire;
  assign TLB_1_or29 = OptimizationBarrier_28_metaAssert_wire | TLB_1_or60;
  assign TLB_1_or62 = OptimizationBarrier_17_metaAssert_wire | OptimizationBarrier_35_metaAssert_wire;
  assign TLB_1_or30 = OptimizationBarrier_23_metaAssert_wire | TLB_1_or62;
  assign TLB_1_or14 = TLB_1_or29 | TLB_1_or30;
  assign TLB_1_or6 = TLB_1_or13 | TLB_1_or14;
  assign TLB_1_or2 = TLB_1_or5 | TLB_1_or6;
  assign TLB_1_or0 = TLB_1_or1 | TLB_1_or2;
  assign metaAssert = TLB_1_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_tag = _RAND_0[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_data_0 = _RAND_1[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_data_1 = _RAND_2[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_data_2 = _RAND_3[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_data_3 = _RAND_4[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_valid_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_valid_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_valid_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_valid_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_1_tag = _RAND_9[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_1_data_0 = _RAND_10[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_1_data_1 = _RAND_11[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_1_data_2 = _RAND_12[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_1_data_3 = _RAND_13[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_1_valid_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_1_valid_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_1_valid_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_1_valid_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sectored_entries_2_tag = _RAND_18[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  sectored_entries_2_data_0 = _RAND_19[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  sectored_entries_2_data_1 = _RAND_20[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  sectored_entries_2_data_2 = _RAND_21[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  sectored_entries_2_data_3 = _RAND_22[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sectored_entries_2_valid_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sectored_entries_2_valid_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sectored_entries_2_valid_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sectored_entries_2_valid_3 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sectored_entries_3_tag = _RAND_27[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  sectored_entries_3_data_0 = _RAND_28[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  sectored_entries_3_data_1 = _RAND_29[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  sectored_entries_3_data_2 = _RAND_30[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  sectored_entries_3_data_3 = _RAND_31[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sectored_entries_3_valid_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sectored_entries_3_valid_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  sectored_entries_3_valid_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  sectored_entries_3_valid_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sectored_entries_4_tag = _RAND_36[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  sectored_entries_4_data_0 = _RAND_37[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  sectored_entries_4_data_1 = _RAND_38[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  sectored_entries_4_data_2 = _RAND_39[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  sectored_entries_4_data_3 = _RAND_40[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  sectored_entries_4_valid_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  sectored_entries_4_valid_1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  sectored_entries_4_valid_2 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  sectored_entries_4_valid_3 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  sectored_entries_5_tag = _RAND_45[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  sectored_entries_5_data_0 = _RAND_46[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  sectored_entries_5_data_1 = _RAND_47[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  sectored_entries_5_data_2 = _RAND_48[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  sectored_entries_5_data_3 = _RAND_49[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  sectored_entries_5_valid_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  sectored_entries_5_valid_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  sectored_entries_5_valid_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  sectored_entries_5_valid_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  sectored_entries_6_tag = _RAND_54[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  sectored_entries_6_data_0 = _RAND_55[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  sectored_entries_6_data_1 = _RAND_56[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  sectored_entries_6_data_2 = _RAND_57[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  sectored_entries_6_data_3 = _RAND_58[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  sectored_entries_6_valid_0 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  sectored_entries_6_valid_1 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  sectored_entries_6_valid_2 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  sectored_entries_6_valid_3 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  sectored_entries_7_tag = _RAND_63[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{`RANDOM}};
  sectored_entries_7_data_0 = _RAND_64[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  sectored_entries_7_data_1 = _RAND_65[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  sectored_entries_7_data_2 = _RAND_66[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  sectored_entries_7_data_3 = _RAND_67[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  sectored_entries_7_valid_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  sectored_entries_7_valid_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  sectored_entries_7_valid_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  sectored_entries_7_valid_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  superpage_entries_0_level = _RAND_72[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_73[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_74[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  superpage_entries_1_level = _RAND_76[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_77[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_78[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  superpage_entries_2_level = _RAND_80[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_81[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_82[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  superpage_entries_3_level = _RAND_84[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_85[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_86[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  special_entry_level = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  special_entry_tag = _RAND_89[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_90[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  state = _RAND_92[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  r_refill_tag = _RAND_93[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_94[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_96[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  r_sectored_hit = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_2116 = _RAND_98[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_2117 = _RAND_99[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  TLB_1_state = _RAND_100[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    TLB_1_cov[initvar] = _RAND_101[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  TLB_1_covSum = _RAND_102[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  TLB_1_metaAssert = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      sectored_entries_0_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1147) begin
            sectored_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1147) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1147) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1147) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1147) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2462) begin
          if (sectored_entries_0_data_0[0]) begin
            sectored_entries_0_valid_0 <= 1'h0;
          end else if (_T_422) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_0_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1147) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_valid_0 <= _GEN_85;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_0 <= _GEN_85;
                  end
                end
              end
            end
          end
        end else if (_T_422) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_0_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_0 <= _GEN_85;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1147) begin
                if (invalidate_refill) begin
                  sectored_entries_0_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_valid_0 <= _GEN_85;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_0 <= _GEN_685;
      end
    end else begin
      sectored_entries_0_valid_0 <= _GEN_505;
    end
    if (metaReset) begin
      sectored_entries_0_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_0_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2462) begin
          if (sectored_entries_0_data_1[0]) begin
            sectored_entries_0_valid_1 <= 1'h0;
          end else if (_T_422) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_0_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1147) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_valid_1 <= _GEN_86;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_1 <= _GEN_86;
                  end
                end
              end
            end
          end
        end else if (_T_422) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_0_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_1 <= _GEN_86;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1147) begin
                if (invalidate_refill) begin
                  sectored_entries_0_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_valid_1 <= _GEN_86;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_1 <= _GEN_686;
      end
    end else begin
      sectored_entries_0_valid_1 <= _GEN_506;
    end
    if (metaReset) begin
      sectored_entries_0_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_0_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2462) begin
          if (sectored_entries_0_data_2[0]) begin
            sectored_entries_0_valid_2 <= 1'h0;
          end else if (_T_422) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_0_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1147) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_valid_2 <= _GEN_87;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_2 <= _GEN_87;
                  end
                end
              end
            end
          end
        end else if (_T_422) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_0_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_2 <= _GEN_87;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1147) begin
                if (invalidate_refill) begin
                  sectored_entries_0_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_valid_2 <= _GEN_87;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_2 <= _GEN_687;
      end
    end else begin
      sectored_entries_0_valid_2 <= _GEN_507;
    end
    if (metaReset) begin
      sectored_entries_0_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_0_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2462) begin
          if (sectored_entries_0_data_3[0]) begin
            sectored_entries_0_valid_3 <= 1'h0;
          end else if (_T_422) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_0_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1147) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_valid_3 <= _GEN_88;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_3 <= _GEN_88;
                  end
                end
              end
            end
          end
        end else if (_T_422) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_0_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1147) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_valid_3 <= _GEN_88;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1147) begin
                if (invalidate_refill) begin
                  sectored_entries_0_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_valid_3 <= _GEN_88;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_3 <= _GEN_688;
      end
    end else begin
      sectored_entries_0_valid_3 <= _GEN_508;
    end
    if (metaReset) begin
      sectored_entries_1_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1165) begin
            sectored_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1165) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1165) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1165) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1165) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2617) begin
          if (sectored_entries_1_data_0[0]) begin
            sectored_entries_1_valid_0 <= 1'h0;
          end else if (_T_428) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_1_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1165) begin
                    if (invalidate_refill) begin
                      sectored_entries_1_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_1_valid_0 <= _GEN_111;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_0 <= _GEN_111;
                  end
                end
              end
            end
          end
        end else if (_T_428) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_1_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_0 <= _GEN_111;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1165) begin
                if (invalidate_refill) begin
                  sectored_entries_1_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_1_valid_0 <= _GEN_111;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_0 <= _GEN_713;
      end
    end else begin
      sectored_entries_1_valid_0 <= _GEN_515;
    end
    if (metaReset) begin
      sectored_entries_1_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_1_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2617) begin
          if (sectored_entries_1_data_1[0]) begin
            sectored_entries_1_valid_1 <= 1'h0;
          end else if (_T_428) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_1_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1165) begin
                    if (invalidate_refill) begin
                      sectored_entries_1_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_1_valid_1 <= _GEN_112;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_1 <= _GEN_112;
                  end
                end
              end
            end
          end
        end else if (_T_428) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_1_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_1 <= _GEN_112;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1165) begin
                if (invalidate_refill) begin
                  sectored_entries_1_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_1_valid_1 <= _GEN_112;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_1 <= _GEN_714;
      end
    end else begin
      sectored_entries_1_valid_1 <= _GEN_516;
    end
    if (metaReset) begin
      sectored_entries_1_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_1_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2617) begin
          if (sectored_entries_1_data_2[0]) begin
            sectored_entries_1_valid_2 <= 1'h0;
          end else if (_T_428) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_1_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1165) begin
                    if (invalidate_refill) begin
                      sectored_entries_1_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_1_valid_2 <= _GEN_113;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_2 <= _GEN_113;
                  end
                end
              end
            end
          end
        end else if (_T_428) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_1_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_2 <= _GEN_113;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1165) begin
                if (invalidate_refill) begin
                  sectored_entries_1_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_1_valid_2 <= _GEN_113;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_2 <= _GEN_715;
      end
    end else begin
      sectored_entries_1_valid_2 <= _GEN_517;
    end
    if (metaReset) begin
      sectored_entries_1_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_1_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2617) begin
          if (sectored_entries_1_data_3[0]) begin
            sectored_entries_1_valid_3 <= 1'h0;
          end else if (_T_428) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_1_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1165) begin
                    if (invalidate_refill) begin
                      sectored_entries_1_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_1_valid_3 <= _GEN_114;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_3 <= _GEN_114;
                  end
                end
              end
            end
          end
        end else if (_T_428) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_1_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1165) begin
                  if (invalidate_refill) begin
                    sectored_entries_1_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_1_valid_3 <= _GEN_114;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1165) begin
                if (invalidate_refill) begin
                  sectored_entries_1_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_1_valid_3 <= _GEN_114;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_3 <= _GEN_716;
      end
    end else begin
      sectored_entries_1_valid_3 <= _GEN_518;
    end
    if (metaReset) begin
      sectored_entries_2_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1183) begin
            sectored_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1183) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1183) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1183) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1183) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2772) begin
          if (sectored_entries_2_data_0[0]) begin
            sectored_entries_2_valid_0 <= 1'h0;
          end else if (_T_434) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_2_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1183) begin
                    if (invalidate_refill) begin
                      sectored_entries_2_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_2_valid_0 <= _GEN_137;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_0 <= _GEN_137;
                  end
                end
              end
            end
          end
        end else if (_T_434) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_2_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_0 <= _GEN_137;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1183) begin
                if (invalidate_refill) begin
                  sectored_entries_2_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_2_valid_0 <= _GEN_137;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_0 <= _GEN_741;
      end
    end else begin
      sectored_entries_2_valid_0 <= _GEN_525;
    end
    if (metaReset) begin
      sectored_entries_2_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_2_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2772) begin
          if (sectored_entries_2_data_1[0]) begin
            sectored_entries_2_valid_1 <= 1'h0;
          end else if (_T_434) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_2_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1183) begin
                    if (invalidate_refill) begin
                      sectored_entries_2_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_2_valid_1 <= _GEN_138;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_1 <= _GEN_138;
                  end
                end
              end
            end
          end
        end else if (_T_434) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_2_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_1 <= _GEN_138;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1183) begin
                if (invalidate_refill) begin
                  sectored_entries_2_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_2_valid_1 <= _GEN_138;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_1 <= _GEN_742;
      end
    end else begin
      sectored_entries_2_valid_1 <= _GEN_526;
    end
    if (metaReset) begin
      sectored_entries_2_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_2_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2772) begin
          if (sectored_entries_2_data_2[0]) begin
            sectored_entries_2_valid_2 <= 1'h0;
          end else if (_T_434) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_2_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1183) begin
                    if (invalidate_refill) begin
                      sectored_entries_2_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_2_valid_2 <= _GEN_139;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_2 <= _GEN_139;
                  end
                end
              end
            end
          end
        end else if (_T_434) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_2_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_2 <= _GEN_139;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1183) begin
                if (invalidate_refill) begin
                  sectored_entries_2_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_2_valid_2 <= _GEN_139;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_2 <= _GEN_743;
      end
    end else begin
      sectored_entries_2_valid_2 <= _GEN_527;
    end
    if (metaReset) begin
      sectored_entries_2_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_2_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2772) begin
          if (sectored_entries_2_data_3[0]) begin
            sectored_entries_2_valid_3 <= 1'h0;
          end else if (_T_434) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_2_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1183) begin
                    if (invalidate_refill) begin
                      sectored_entries_2_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_2_valid_3 <= _GEN_140;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_3 <= _GEN_140;
                  end
                end
              end
            end
          end
        end else if (_T_434) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_2_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1183) begin
                  if (invalidate_refill) begin
                    sectored_entries_2_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_2_valid_3 <= _GEN_140;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1183) begin
                if (invalidate_refill) begin
                  sectored_entries_2_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_2_valid_3 <= _GEN_140;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_3 <= _GEN_744;
      end
    end else begin
      sectored_entries_2_valid_3 <= _GEN_528;
    end
    if (metaReset) begin
      sectored_entries_3_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1201) begin
            sectored_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1201) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1201) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1201) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1201) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2927) begin
          if (sectored_entries_3_data_0[0]) begin
            sectored_entries_3_valid_0 <= 1'h0;
          end else if (_T_440) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_3_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1201) begin
                    if (invalidate_refill) begin
                      sectored_entries_3_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_3_valid_0 <= _GEN_163;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_0 <= _GEN_163;
                  end
                end
              end
            end
          end
        end else if (_T_440) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_3_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_0 <= _GEN_163;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1201) begin
                if (invalidate_refill) begin
                  sectored_entries_3_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_3_valid_0 <= _GEN_163;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_0 <= _GEN_769;
      end
    end else begin
      sectored_entries_3_valid_0 <= _GEN_535;
    end
    if (metaReset) begin
      sectored_entries_3_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_3_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2927) begin
          if (sectored_entries_3_data_1[0]) begin
            sectored_entries_3_valid_1 <= 1'h0;
          end else if (_T_440) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_3_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1201) begin
                    if (invalidate_refill) begin
                      sectored_entries_3_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_3_valid_1 <= _GEN_164;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_1 <= _GEN_164;
                  end
                end
              end
            end
          end
        end else if (_T_440) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_3_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_1 <= _GEN_164;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1201) begin
                if (invalidate_refill) begin
                  sectored_entries_3_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_3_valid_1 <= _GEN_164;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_1 <= _GEN_770;
      end
    end else begin
      sectored_entries_3_valid_1 <= _GEN_536;
    end
    if (metaReset) begin
      sectored_entries_3_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_3_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2927) begin
          if (sectored_entries_3_data_2[0]) begin
            sectored_entries_3_valid_2 <= 1'h0;
          end else if (_T_440) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_3_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1201) begin
                    if (invalidate_refill) begin
                      sectored_entries_3_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_3_valid_2 <= _GEN_165;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_2 <= _GEN_165;
                  end
                end
              end
            end
          end
        end else if (_T_440) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_3_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_2 <= _GEN_165;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1201) begin
                if (invalidate_refill) begin
                  sectored_entries_3_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_3_valid_2 <= _GEN_165;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_2 <= _GEN_771;
      end
    end else begin
      sectored_entries_3_valid_2 <= _GEN_537;
    end
    if (metaReset) begin
      sectored_entries_3_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_3_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2927) begin
          if (sectored_entries_3_data_3[0]) begin
            sectored_entries_3_valid_3 <= 1'h0;
          end else if (_T_440) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_3_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1201) begin
                    if (invalidate_refill) begin
                      sectored_entries_3_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_3_valid_3 <= _GEN_166;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_3 <= _GEN_166;
                  end
                end
              end
            end
          end
        end else if (_T_440) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_3_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1201) begin
                  if (invalidate_refill) begin
                    sectored_entries_3_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_3_valid_3 <= _GEN_166;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1201) begin
                if (invalidate_refill) begin
                  sectored_entries_3_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_3_valid_3 <= _GEN_166;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_3 <= _GEN_772;
      end
    end else begin
      sectored_entries_3_valid_3 <= _GEN_538;
    end
    if (metaReset) begin
      sectored_entries_4_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1219) begin
            sectored_entries_4_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1219) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1219) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1219) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1219) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_4_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3082) begin
          if (sectored_entries_4_data_0[0]) begin
            sectored_entries_4_valid_0 <= 1'h0;
          end else if (_T_446) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_4_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1219) begin
                    if (invalidate_refill) begin
                      sectored_entries_4_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_4_valid_0 <= _GEN_189;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_0 <= _GEN_189;
                  end
                end
              end
            end
          end
        end else if (_T_446) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_4_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_0 <= _GEN_189;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1219) begin
                if (invalidate_refill) begin
                  sectored_entries_4_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_4_valid_0 <= _GEN_189;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_0 <= _GEN_797;
      end
    end else begin
      sectored_entries_4_valid_0 <= _GEN_545;
    end
    if (metaReset) begin
      sectored_entries_4_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_4_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3082) begin
          if (sectored_entries_4_data_1[0]) begin
            sectored_entries_4_valid_1 <= 1'h0;
          end else if (_T_446) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_4_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1219) begin
                    if (invalidate_refill) begin
                      sectored_entries_4_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_4_valid_1 <= _GEN_190;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_1 <= _GEN_190;
                  end
                end
              end
            end
          end
        end else if (_T_446) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_4_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_1 <= _GEN_190;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1219) begin
                if (invalidate_refill) begin
                  sectored_entries_4_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_4_valid_1 <= _GEN_190;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_1 <= _GEN_798;
      end
    end else begin
      sectored_entries_4_valid_1 <= _GEN_546;
    end
    if (metaReset) begin
      sectored_entries_4_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_4_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3082) begin
          if (sectored_entries_4_data_2[0]) begin
            sectored_entries_4_valid_2 <= 1'h0;
          end else if (_T_446) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_4_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1219) begin
                    if (invalidate_refill) begin
                      sectored_entries_4_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_4_valid_2 <= _GEN_191;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_2 <= _GEN_191;
                  end
                end
              end
            end
          end
        end else if (_T_446) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_4_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_2 <= _GEN_191;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1219) begin
                if (invalidate_refill) begin
                  sectored_entries_4_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_4_valid_2 <= _GEN_191;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_2 <= _GEN_799;
      end
    end else begin
      sectored_entries_4_valid_2 <= _GEN_547;
    end
    if (metaReset) begin
      sectored_entries_4_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_4_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3082) begin
          if (sectored_entries_4_data_3[0]) begin
            sectored_entries_4_valid_3 <= 1'h0;
          end else if (_T_446) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_4_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1219) begin
                    if (invalidate_refill) begin
                      sectored_entries_4_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_4_valid_3 <= _GEN_192;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_3 <= _GEN_192;
                  end
                end
              end
            end
          end
        end else if (_T_446) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_4_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1219) begin
                  if (invalidate_refill) begin
                    sectored_entries_4_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_4_valid_3 <= _GEN_192;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1219) begin
                if (invalidate_refill) begin
                  sectored_entries_4_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_4_valid_3 <= _GEN_192;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_3 <= _GEN_800;
      end
    end else begin
      sectored_entries_4_valid_3 <= _GEN_548;
    end
    if (metaReset) begin
      sectored_entries_5_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1237) begin
            sectored_entries_5_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1237) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1237) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1237) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1237) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_5_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3237) begin
          if (sectored_entries_5_data_0[0]) begin
            sectored_entries_5_valid_0 <= 1'h0;
          end else if (_T_452) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_5_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1237) begin
                    if (invalidate_refill) begin
                      sectored_entries_5_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_5_valid_0 <= _GEN_215;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_0 <= _GEN_215;
                  end
                end
              end
            end
          end
        end else if (_T_452) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_5_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_0 <= _GEN_215;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1237) begin
                if (invalidate_refill) begin
                  sectored_entries_5_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_5_valid_0 <= _GEN_215;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_0 <= _GEN_825;
      end
    end else begin
      sectored_entries_5_valid_0 <= _GEN_555;
    end
    if (metaReset) begin
      sectored_entries_5_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_5_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3237) begin
          if (sectored_entries_5_data_1[0]) begin
            sectored_entries_5_valid_1 <= 1'h0;
          end else if (_T_452) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_5_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1237) begin
                    if (invalidate_refill) begin
                      sectored_entries_5_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_5_valid_1 <= _GEN_216;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_1 <= _GEN_216;
                  end
                end
              end
            end
          end
        end else if (_T_452) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_5_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_1 <= _GEN_216;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1237) begin
                if (invalidate_refill) begin
                  sectored_entries_5_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_5_valid_1 <= _GEN_216;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_1 <= _GEN_826;
      end
    end else begin
      sectored_entries_5_valid_1 <= _GEN_556;
    end
    if (metaReset) begin
      sectored_entries_5_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_5_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3237) begin
          if (sectored_entries_5_data_2[0]) begin
            sectored_entries_5_valid_2 <= 1'h0;
          end else if (_T_452) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_5_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1237) begin
                    if (invalidate_refill) begin
                      sectored_entries_5_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_5_valid_2 <= _GEN_217;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_2 <= _GEN_217;
                  end
                end
              end
            end
          end
        end else if (_T_452) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_5_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_2 <= _GEN_217;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1237) begin
                if (invalidate_refill) begin
                  sectored_entries_5_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_5_valid_2 <= _GEN_217;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_2 <= _GEN_827;
      end
    end else begin
      sectored_entries_5_valid_2 <= _GEN_557;
    end
    if (metaReset) begin
      sectored_entries_5_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_5_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3237) begin
          if (sectored_entries_5_data_3[0]) begin
            sectored_entries_5_valid_3 <= 1'h0;
          end else if (_T_452) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_5_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1237) begin
                    if (invalidate_refill) begin
                      sectored_entries_5_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_5_valid_3 <= _GEN_218;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_3 <= _GEN_218;
                  end
                end
              end
            end
          end
        end else if (_T_452) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_5_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1237) begin
                  if (invalidate_refill) begin
                    sectored_entries_5_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_5_valid_3 <= _GEN_218;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1237) begin
                if (invalidate_refill) begin
                  sectored_entries_5_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_5_valid_3 <= _GEN_218;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_3 <= _GEN_828;
      end
    end else begin
      sectored_entries_5_valid_3 <= _GEN_558;
    end
    if (metaReset) begin
      sectored_entries_6_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1255) begin
            sectored_entries_6_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1255) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1255) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1255) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1255) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_6_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3392) begin
          if (sectored_entries_6_data_0[0]) begin
            sectored_entries_6_valid_0 <= 1'h0;
          end else if (_T_458) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_6_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1255) begin
                    if (invalidate_refill) begin
                      sectored_entries_6_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_6_valid_0 <= _GEN_241;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_0 <= _GEN_241;
                  end
                end
              end
            end
          end
        end else if (_T_458) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_6_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_0 <= _GEN_241;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1255) begin
                if (invalidate_refill) begin
                  sectored_entries_6_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_6_valid_0 <= _GEN_241;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_0 <= _GEN_853;
      end
    end else begin
      sectored_entries_6_valid_0 <= _GEN_565;
    end
    if (metaReset) begin
      sectored_entries_6_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_6_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3392) begin
          if (sectored_entries_6_data_1[0]) begin
            sectored_entries_6_valid_1 <= 1'h0;
          end else if (_T_458) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_6_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1255) begin
                    if (invalidate_refill) begin
                      sectored_entries_6_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_6_valid_1 <= _GEN_242;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_1 <= _GEN_242;
                  end
                end
              end
            end
          end
        end else if (_T_458) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_6_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_1 <= _GEN_242;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1255) begin
                if (invalidate_refill) begin
                  sectored_entries_6_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_6_valid_1 <= _GEN_242;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_1 <= _GEN_854;
      end
    end else begin
      sectored_entries_6_valid_1 <= _GEN_566;
    end
    if (metaReset) begin
      sectored_entries_6_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_6_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3392) begin
          if (sectored_entries_6_data_2[0]) begin
            sectored_entries_6_valid_2 <= 1'h0;
          end else if (_T_458) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_6_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1255) begin
                    if (invalidate_refill) begin
                      sectored_entries_6_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_6_valid_2 <= _GEN_243;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_2 <= _GEN_243;
                  end
                end
              end
            end
          end
        end else if (_T_458) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_6_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_2 <= _GEN_243;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1255) begin
                if (invalidate_refill) begin
                  sectored_entries_6_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_6_valid_2 <= _GEN_243;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_2 <= _GEN_855;
      end
    end else begin
      sectored_entries_6_valid_2 <= _GEN_567;
    end
    if (metaReset) begin
      sectored_entries_6_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_6_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3392) begin
          if (sectored_entries_6_data_3[0]) begin
            sectored_entries_6_valid_3 <= 1'h0;
          end else if (_T_458) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_6_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1255) begin
                    if (invalidate_refill) begin
                      sectored_entries_6_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_6_valid_3 <= _GEN_244;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_3 <= _GEN_244;
                  end
                end
              end
            end
          end
        end else if (_T_458) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_6_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1255) begin
                  if (invalidate_refill) begin
                    sectored_entries_6_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_6_valid_3 <= _GEN_244;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1255) begin
                if (invalidate_refill) begin
                  sectored_entries_6_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_6_valid_3 <= _GEN_244;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_3 <= _GEN_856;
      end
    end else begin
      sectored_entries_6_valid_3 <= _GEN_568;
    end
    if (metaReset) begin
      sectored_entries_7_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1273) begin
            sectored_entries_7_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1273) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_0 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1273) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_1 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1273) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_2 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1077)) begin
          if (_T_1273) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_3 <= _T_1076;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_7_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3547) begin
          if (sectored_entries_7_data_0[0]) begin
            sectored_entries_7_valid_0 <= 1'h0;
          end else if (_T_464) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_7_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1273) begin
                    if (invalidate_refill) begin
                      sectored_entries_7_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_7_valid_0 <= _GEN_267;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_0 <= _GEN_267;
                  end
                end
              end
            end
          end
        end else if (_T_464) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_7_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_0 <= _GEN_267;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1273) begin
                if (invalidate_refill) begin
                  sectored_entries_7_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_7_valid_0 <= _GEN_267;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_0 <= _GEN_881;
      end
    end else begin
      sectored_entries_7_valid_0 <= _GEN_575;
    end
    if (metaReset) begin
      sectored_entries_7_valid_1 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_7_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3547) begin
          if (sectored_entries_7_data_1[0]) begin
            sectored_entries_7_valid_1 <= 1'h0;
          end else if (_T_464) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_7_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1273) begin
                    if (invalidate_refill) begin
                      sectored_entries_7_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_7_valid_1 <= _GEN_268;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_1 <= _GEN_268;
                  end
                end
              end
            end
          end
        end else if (_T_464) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_7_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_1 <= _GEN_268;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1273) begin
                if (invalidate_refill) begin
                  sectored_entries_7_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_7_valid_1 <= _GEN_268;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_1 <= _GEN_882;
      end
    end else begin
      sectored_entries_7_valid_1 <= _GEN_576;
    end
    if (metaReset) begin
      sectored_entries_7_valid_2 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_7_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3547) begin
          if (sectored_entries_7_data_2[0]) begin
            sectored_entries_7_valid_2 <= 1'h0;
          end else if (_T_464) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_7_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1273) begin
                    if (invalidate_refill) begin
                      sectored_entries_7_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_7_valid_2 <= _GEN_269;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_2 <= _GEN_269;
                  end
                end
              end
            end
          end
        end else if (_T_464) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_7_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_2 <= _GEN_269;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1273) begin
                if (invalidate_refill) begin
                  sectored_entries_7_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_7_valid_2 <= _GEN_269;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_2 <= _GEN_883;
      end
    end else begin
      sectored_entries_7_valid_2 <= _GEN_577;
    end
    if (metaReset) begin
      sectored_entries_7_valid_3 <= 1'h0;
    end else if (_T_3897) begin
      sectored_entries_7_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3547) begin
          if (sectored_entries_7_data_3[0]) begin
            sectored_entries_7_valid_3 <= 1'h0;
          end else if (_T_464) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_7_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1077)) begin
                  if (_T_1273) begin
                    if (invalidate_refill) begin
                      sectored_entries_7_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_7_valid_3 <= _GEN_270;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_3 <= _GEN_270;
                  end
                end
              end
            end
          end
        end else if (_T_464) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_7_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1077)) begin
                if (_T_1273) begin
                  if (invalidate_refill) begin
                    sectored_entries_7_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_7_valid_3 <= _GEN_270;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1077)) begin
              if (_T_1273) begin
                if (invalidate_refill) begin
                  sectored_entries_7_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_7_valid_3 <= _GEN_270;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_3 <= _GEN_884;
      end
    end else begin
      sectored_entries_7_valid_3 <= _GEN_578;
    end
    if (metaReset) begin
      superpage_entries_0_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1078) begin
            superpage_entries_0_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1078) begin
            superpage_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1078) begin
            superpage_entries_0_data_0 <= _T_1076;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_0) begin
          superpage_entries_0_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1077) begin
              if (_T_1078) begin
                if (invalidate_refill) begin
                  superpage_entries_0_valid_0 <= 1'h0;
                end else begin
                  superpage_entries_0_valid_0 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        superpage_entries_0_valid_0 <= _GEN_891;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1078) begin
            if (invalidate_refill) begin
              superpage_entries_0_valid_0 <= 1'h0;
            end else begin
              superpage_entries_0_valid_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1095) begin
            superpage_entries_1_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1095) begin
            superpage_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1095) begin
            superpage_entries_1_data_0 <= _T_1076;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_1) begin
          superpage_entries_1_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1077) begin
              if (_T_1095) begin
                if (invalidate_refill) begin
                  superpage_entries_1_valid_0 <= 1'h0;
                end else begin
                  superpage_entries_1_valid_0 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        superpage_entries_1_valid_0 <= _GEN_895;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1095) begin
            if (invalidate_refill) begin
              superpage_entries_1_valid_0 <= 1'h0;
            end else begin
              superpage_entries_1_valid_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1112) begin
            superpage_entries_2_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1112) begin
            superpage_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1112) begin
            superpage_entries_2_data_0 <= _T_1076;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_2) begin
          superpage_entries_2_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1077) begin
              if (_T_1112) begin
                superpage_entries_2_valid_0 <= _GEN_64;
              end
            end
          end
        end
      end else begin
        superpage_entries_2_valid_0 <= _GEN_899;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1112) begin
            superpage_entries_2_valid_0 <= _GEN_64;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1129) begin
            superpage_entries_3_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1129) begin
            superpage_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1129) begin
            superpage_entries_3_data_0 <= _T_1076;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_3) begin
          superpage_entries_3_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1077) begin
              if (_T_1129) begin
                superpage_entries_3_valid_0 <= _GEN_64;
              end
            end
          end
        end
      end else begin
        superpage_entries_3_valid_0 <= _GEN_903;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1077) begin
          if (_T_1129) begin
            superpage_entries_3_valid_0 <= _GEN_64;
          end
        end
      end
    end
    if (metaReset) begin
      special_entry_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_level <= io_ptw_resp_bits_level;
      end
    end
    if (metaReset) begin
      special_entry_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_tag <= r_refill_tag;
      end
    end
    if (metaReset) begin
      special_entry_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_data_0 <= _T_1076;
      end
    end
    if (metaReset) begin
      special_entry_valid_0 <= 1'h0;
    end else if (_T_3897) begin
      special_entry_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_689) begin
          special_entry_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (~io_ptw_resp_bits_homogeneous) begin
            special_entry_valid_0 <= _GEN_64;
          end
        end
      end else begin
        special_entry_valid_0 <= _GEN_907;
      end
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_valid_0 <= _GEN_64;
      end
    end
    if (metaReset) begin
      state <= 2'h0;
    end else if (reset) begin
      state <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if (_T_2448) begin
      state <= 2'h3;
    end else if (_T_4) begin
      if (io_kill) begin
        state <= 2'h0;
      end else if (io_ptw_req_ready) begin
        if (io_sfence_valid) begin
          state <= 2'h3;
        end else begin
          state <= 2'h2;
        end
      end else if (io_sfence_valid) begin
        state <= 2'h0;
      end else if (_T_2331) begin
        state <= 2'h1;
      end
    end else if (_T_2331) begin
      state <= 2'h1;
    end
    if (metaReset) begin
      r_refill_tag <= 27'h0;
    end else if (_T_2331) begin
      r_refill_tag <= vpn;
    end
    if (metaReset) begin
      r_superpage_repl_addr <= 2'h0;
    end else if (_T_2331) begin
      if (_T_2342) begin
        r_superpage_repl_addr <= _T_2338;
      end else if (_T_2344) begin
        r_superpage_repl_addr <= 2'h0;
      end else if (_T_2345) begin
        r_superpage_repl_addr <= 2'h1;
      end else if (_T_2346) begin
        r_superpage_repl_addr <= 2'h2;
      end else begin
        r_superpage_repl_addr <= 2'h3;
      end
    end
    if (metaReset) begin
      r_sectored_repl_addr <= 3'h0;
    end else if (_T_2331) begin
      if (_T_2402) begin
        r_sectored_repl_addr <= _T_2370;
      end else if (_T_2404) begin
        r_sectored_repl_addr <= 3'h0;
      end else if (_T_2405) begin
        r_sectored_repl_addr <= 3'h1;
      end else if (_T_2406) begin
        r_sectored_repl_addr <= 3'h2;
      end else if (_T_2407) begin
        r_sectored_repl_addr <= 3'h3;
      end else if (_T_2408) begin
        r_sectored_repl_addr <= 3'h4;
      end else if (_T_2409) begin
        r_sectored_repl_addr <= 3'h5;
      end else if (_T_2410) begin
        r_sectored_repl_addr <= 3'h6;
      end else begin
        r_sectored_repl_addr <= 3'h7;
      end
    end
    if (metaReset) begin
      r_sectored_hit_addr <= 3'h0;
    end else if (_T_2331) begin
      r_sectored_hit_addr <= _T_2143;
    end
    if (metaReset) begin
      r_sectored_hit <= 1'h0;
    end else if (_T_2331) begin
      r_sectored_hit <= _T_2125;
    end
    if (metaReset) begin
      _T_2116 <= 7'h0;
    end else if (_T_2118) begin
      if (_T_2125) begin
        _T_2116 <= _T_2182;
      end
    end
    if (metaReset) begin
      _T_2117 <= 3'h0;
    end else if (_T_2118) begin
      if (_T_2185) begin
        _T_2117 <= _T_2209;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & ~_T_2454) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:381 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"); // @[TLB.scala 381:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_sfence_valid & ~_T_2454) begin
          $fatal; // @[TLB.scala 381:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    TLB_1_state <= TLB_1_xor0;
    if (!(TLB_1_cov_read_data)) begin
      TLB_1_covSum <= TLB_1_covSum + 1'h1;
    end
    if (metaReset) begin
      TLB_1_metaAssert <= 1'h0;
    end else begin
      TLB_1_metaAssert <= TLB_1_metaAssert | TLB_1_or0;
    end
  end
  always @(posedge clock) begin
    if(TLB_1_cov_write_en & TLB_1_cov_write_mask) begin
      TLB_1_cov[TLB_1_cov_write_addr] <= TLB_1_cov_write_data; // @[Coverage map for TLB_1]
    end
  end
endmodule
module BTB(
  input         clock,
  input         reset,
  input  [38:0] io_req_bits_addr,
  output        io_resp_valid,
  output        io_resp_bits_taken,
  output        io_resp_bits_bridx,
  output [38:0] io_resp_bits_target,
  output [4:0]  io_resp_bits_entry,
  output [7:0]  io_resp_bits_bht_history,
  output        io_resp_bits_bht_value,
  input         io_btb_update_valid,
  input  [4:0]  io_btb_update_bits_prediction_entry,
  input  [38:0] io_btb_update_bits_pc,
  input         io_btb_update_bits_isValid,
  input  [38:0] io_btb_update_bits_br_pc,
  input  [1:0]  io_btb_update_bits_cfiType,
  input         io_bht_update_valid,
  input  [7:0]  io_bht_update_bits_prediction_history,
  input  [38:0] io_bht_update_bits_pc,
  input         io_bht_update_bits_branch,
  input         io_bht_update_bits_taken,
  input         io_bht_update_bits_mispredict,
  input         io_bht_advance_valid,
  input         io_bht_advance_bits_bht_value,
  input         io_ras_update_valid,
  input  [1:0]  io_ras_update_bits_cfiType,
  input  [38:0] io_ras_update_bits_returnAddr,
  output        io_ras_head_valid,
  output [38:0] io_ras_head_bits,
  input         io_flush,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  _T_1037 [0:511]; // @[BTB.scala 113:26]
  reg [31:0] _RAND_0;
  wire  _T_1037__T_1106_data; // @[BTB.scala 113:26]
  wire [8:0] _T_1037__T_1106_addr; // @[BTB.scala 113:26]
  wire  _T_1037__T_1119_data; // @[BTB.scala 113:26]
  wire [8:0] _T_1037__T_1119_addr; // @[BTB.scala 113:26]
  wire  _T_1037__T_1119_mask; // @[BTB.scala 113:26]
  wire  _T_1037__T_1119_en; // @[BTB.scala 113:26]
  reg [12:0] idxs_0; // @[BTB.scala 188:17]
  reg [31:0] _RAND_1;
  reg [12:0] idxs_1; // @[BTB.scala 188:17]
  reg [31:0] _RAND_2;
  reg [12:0] idxs_2; // @[BTB.scala 188:17]
  reg [31:0] _RAND_3;
  reg [12:0] idxs_3; // @[BTB.scala 188:17]
  reg [31:0] _RAND_4;
  reg [12:0] idxs_4; // @[BTB.scala 188:17]
  reg [31:0] _RAND_5;
  reg [12:0] idxs_5; // @[BTB.scala 188:17]
  reg [31:0] _RAND_6;
  reg [12:0] idxs_6; // @[BTB.scala 188:17]
  reg [31:0] _RAND_7;
  reg [12:0] idxs_7; // @[BTB.scala 188:17]
  reg [31:0] _RAND_8;
  reg [12:0] idxs_8; // @[BTB.scala 188:17]
  reg [31:0] _RAND_9;
  reg [12:0] idxs_9; // @[BTB.scala 188:17]
  reg [31:0] _RAND_10;
  reg [12:0] idxs_10; // @[BTB.scala 188:17]
  reg [31:0] _RAND_11;
  reg [12:0] idxs_11; // @[BTB.scala 188:17]
  reg [31:0] _RAND_12;
  reg [12:0] idxs_12; // @[BTB.scala 188:17]
  reg [31:0] _RAND_13;
  reg [12:0] idxs_13; // @[BTB.scala 188:17]
  reg [31:0] _RAND_14;
  reg [12:0] idxs_14; // @[BTB.scala 188:17]
  reg [31:0] _RAND_15;
  reg [12:0] idxs_15; // @[BTB.scala 188:17]
  reg [31:0] _RAND_16;
  reg [12:0] idxs_16; // @[BTB.scala 188:17]
  reg [31:0] _RAND_17;
  reg [12:0] idxs_17; // @[BTB.scala 188:17]
  reg [31:0] _RAND_18;
  reg [12:0] idxs_18; // @[BTB.scala 188:17]
  reg [31:0] _RAND_19;
  reg [12:0] idxs_19; // @[BTB.scala 188:17]
  reg [31:0] _RAND_20;
  reg [12:0] idxs_20; // @[BTB.scala 188:17]
  reg [31:0] _RAND_21;
  reg [12:0] idxs_21; // @[BTB.scala 188:17]
  reg [31:0] _RAND_22;
  reg [12:0] idxs_22; // @[BTB.scala 188:17]
  reg [31:0] _RAND_23;
  reg [12:0] idxs_23; // @[BTB.scala 188:17]
  reg [31:0] _RAND_24;
  reg [12:0] idxs_24; // @[BTB.scala 188:17]
  reg [31:0] _RAND_25;
  reg [12:0] idxs_25; // @[BTB.scala 188:17]
  reg [31:0] _RAND_26;
  reg [12:0] idxs_26; // @[BTB.scala 188:17]
  reg [31:0] _RAND_27;
  reg [12:0] idxs_27; // @[BTB.scala 188:17]
  reg [31:0] _RAND_28;
  reg [2:0] idxPages_0; // @[BTB.scala 189:21]
  reg [31:0] _RAND_29;
  reg [2:0] idxPages_1; // @[BTB.scala 189:21]
  reg [31:0] _RAND_30;
  reg [2:0] idxPages_2; // @[BTB.scala 189:21]
  reg [31:0] _RAND_31;
  reg [2:0] idxPages_3; // @[BTB.scala 189:21]
  reg [31:0] _RAND_32;
  reg [2:0] idxPages_4; // @[BTB.scala 189:21]
  reg [31:0] _RAND_33;
  reg [2:0] idxPages_5; // @[BTB.scala 189:21]
  reg [31:0] _RAND_34;
  reg [2:0] idxPages_6; // @[BTB.scala 189:21]
  reg [31:0] _RAND_35;
  reg [2:0] idxPages_7; // @[BTB.scala 189:21]
  reg [31:0] _RAND_36;
  reg [2:0] idxPages_8; // @[BTB.scala 189:21]
  reg [31:0] _RAND_37;
  reg [2:0] idxPages_9; // @[BTB.scala 189:21]
  reg [31:0] _RAND_38;
  reg [2:0] idxPages_10; // @[BTB.scala 189:21]
  reg [31:0] _RAND_39;
  reg [2:0] idxPages_11; // @[BTB.scala 189:21]
  reg [31:0] _RAND_40;
  reg [2:0] idxPages_12; // @[BTB.scala 189:21]
  reg [31:0] _RAND_41;
  reg [2:0] idxPages_13; // @[BTB.scala 189:21]
  reg [31:0] _RAND_42;
  reg [2:0] idxPages_14; // @[BTB.scala 189:21]
  reg [31:0] _RAND_43;
  reg [2:0] idxPages_15; // @[BTB.scala 189:21]
  reg [31:0] _RAND_44;
  reg [2:0] idxPages_16; // @[BTB.scala 189:21]
  reg [31:0] _RAND_45;
  reg [2:0] idxPages_17; // @[BTB.scala 189:21]
  reg [31:0] _RAND_46;
  reg [2:0] idxPages_18; // @[BTB.scala 189:21]
  reg [31:0] _RAND_47;
  reg [2:0] idxPages_19; // @[BTB.scala 189:21]
  reg [31:0] _RAND_48;
  reg [2:0] idxPages_20; // @[BTB.scala 189:21]
  reg [31:0] _RAND_49;
  reg [2:0] idxPages_21; // @[BTB.scala 189:21]
  reg [31:0] _RAND_50;
  reg [2:0] idxPages_22; // @[BTB.scala 189:21]
  reg [31:0] _RAND_51;
  reg [2:0] idxPages_23; // @[BTB.scala 189:21]
  reg [31:0] _RAND_52;
  reg [2:0] idxPages_24; // @[BTB.scala 189:21]
  reg [31:0] _RAND_53;
  reg [2:0] idxPages_25; // @[BTB.scala 189:21]
  reg [31:0] _RAND_54;
  reg [2:0] idxPages_26; // @[BTB.scala 189:21]
  reg [31:0] _RAND_55;
  reg [2:0] idxPages_27; // @[BTB.scala 189:21]
  reg [31:0] _RAND_56;
  reg [12:0] tgts_0; // @[BTB.scala 190:17]
  reg [31:0] _RAND_57;
  reg [12:0] tgts_1; // @[BTB.scala 190:17]
  reg [31:0] _RAND_58;
  reg [12:0] tgts_2; // @[BTB.scala 190:17]
  reg [31:0] _RAND_59;
  reg [12:0] tgts_3; // @[BTB.scala 190:17]
  reg [31:0] _RAND_60;
  reg [12:0] tgts_4; // @[BTB.scala 190:17]
  reg [31:0] _RAND_61;
  reg [12:0] tgts_5; // @[BTB.scala 190:17]
  reg [31:0] _RAND_62;
  reg [12:0] tgts_6; // @[BTB.scala 190:17]
  reg [31:0] _RAND_63;
  reg [12:0] tgts_7; // @[BTB.scala 190:17]
  reg [31:0] _RAND_64;
  reg [12:0] tgts_8; // @[BTB.scala 190:17]
  reg [31:0] _RAND_65;
  reg [12:0] tgts_9; // @[BTB.scala 190:17]
  reg [31:0] _RAND_66;
  reg [12:0] tgts_10; // @[BTB.scala 190:17]
  reg [31:0] _RAND_67;
  reg [12:0] tgts_11; // @[BTB.scala 190:17]
  reg [31:0] _RAND_68;
  reg [12:0] tgts_12; // @[BTB.scala 190:17]
  reg [31:0] _RAND_69;
  reg [12:0] tgts_13; // @[BTB.scala 190:17]
  reg [31:0] _RAND_70;
  reg [12:0] tgts_14; // @[BTB.scala 190:17]
  reg [31:0] _RAND_71;
  reg [12:0] tgts_15; // @[BTB.scala 190:17]
  reg [31:0] _RAND_72;
  reg [12:0] tgts_16; // @[BTB.scala 190:17]
  reg [31:0] _RAND_73;
  reg [12:0] tgts_17; // @[BTB.scala 190:17]
  reg [31:0] _RAND_74;
  reg [12:0] tgts_18; // @[BTB.scala 190:17]
  reg [31:0] _RAND_75;
  reg [12:0] tgts_19; // @[BTB.scala 190:17]
  reg [31:0] _RAND_76;
  reg [12:0] tgts_20; // @[BTB.scala 190:17]
  reg [31:0] _RAND_77;
  reg [12:0] tgts_21; // @[BTB.scala 190:17]
  reg [31:0] _RAND_78;
  reg [12:0] tgts_22; // @[BTB.scala 190:17]
  reg [31:0] _RAND_79;
  reg [12:0] tgts_23; // @[BTB.scala 190:17]
  reg [31:0] _RAND_80;
  reg [12:0] tgts_24; // @[BTB.scala 190:17]
  reg [31:0] _RAND_81;
  reg [12:0] tgts_25; // @[BTB.scala 190:17]
  reg [31:0] _RAND_82;
  reg [12:0] tgts_26; // @[BTB.scala 190:17]
  reg [31:0] _RAND_83;
  reg [12:0] tgts_27; // @[BTB.scala 190:17]
  reg [31:0] _RAND_84;
  reg [2:0] tgtPages_0; // @[BTB.scala 191:21]
  reg [31:0] _RAND_85;
  reg [2:0] tgtPages_1; // @[BTB.scala 191:21]
  reg [31:0] _RAND_86;
  reg [2:0] tgtPages_2; // @[BTB.scala 191:21]
  reg [31:0] _RAND_87;
  reg [2:0] tgtPages_3; // @[BTB.scala 191:21]
  reg [31:0] _RAND_88;
  reg [2:0] tgtPages_4; // @[BTB.scala 191:21]
  reg [31:0] _RAND_89;
  reg [2:0] tgtPages_5; // @[BTB.scala 191:21]
  reg [31:0] _RAND_90;
  reg [2:0] tgtPages_6; // @[BTB.scala 191:21]
  reg [31:0] _RAND_91;
  reg [2:0] tgtPages_7; // @[BTB.scala 191:21]
  reg [31:0] _RAND_92;
  reg [2:0] tgtPages_8; // @[BTB.scala 191:21]
  reg [31:0] _RAND_93;
  reg [2:0] tgtPages_9; // @[BTB.scala 191:21]
  reg [31:0] _RAND_94;
  reg [2:0] tgtPages_10; // @[BTB.scala 191:21]
  reg [31:0] _RAND_95;
  reg [2:0] tgtPages_11; // @[BTB.scala 191:21]
  reg [31:0] _RAND_96;
  reg [2:0] tgtPages_12; // @[BTB.scala 191:21]
  reg [31:0] _RAND_97;
  reg [2:0] tgtPages_13; // @[BTB.scala 191:21]
  reg [31:0] _RAND_98;
  reg [2:0] tgtPages_14; // @[BTB.scala 191:21]
  reg [31:0] _RAND_99;
  reg [2:0] tgtPages_15; // @[BTB.scala 191:21]
  reg [31:0] _RAND_100;
  reg [2:0] tgtPages_16; // @[BTB.scala 191:21]
  reg [31:0] _RAND_101;
  reg [2:0] tgtPages_17; // @[BTB.scala 191:21]
  reg [31:0] _RAND_102;
  reg [2:0] tgtPages_18; // @[BTB.scala 191:21]
  reg [31:0] _RAND_103;
  reg [2:0] tgtPages_19; // @[BTB.scala 191:21]
  reg [31:0] _RAND_104;
  reg [2:0] tgtPages_20; // @[BTB.scala 191:21]
  reg [31:0] _RAND_105;
  reg [2:0] tgtPages_21; // @[BTB.scala 191:21]
  reg [31:0] _RAND_106;
  reg [2:0] tgtPages_22; // @[BTB.scala 191:21]
  reg [31:0] _RAND_107;
  reg [2:0] tgtPages_23; // @[BTB.scala 191:21]
  reg [31:0] _RAND_108;
  reg [2:0] tgtPages_24; // @[BTB.scala 191:21]
  reg [31:0] _RAND_109;
  reg [2:0] tgtPages_25; // @[BTB.scala 191:21]
  reg [31:0] _RAND_110;
  reg [2:0] tgtPages_26; // @[BTB.scala 191:21]
  reg [31:0] _RAND_111;
  reg [2:0] tgtPages_27; // @[BTB.scala 191:21]
  reg [31:0] _RAND_112;
  reg [24:0] pages_0; // @[BTB.scala 192:18]
  reg [31:0] _RAND_113;
  reg [24:0] pages_1; // @[BTB.scala 192:18]
  reg [31:0] _RAND_114;
  reg [24:0] pages_2; // @[BTB.scala 192:18]
  reg [31:0] _RAND_115;
  reg [24:0] pages_3; // @[BTB.scala 192:18]
  reg [31:0] _RAND_116;
  reg [24:0] pages_4; // @[BTB.scala 192:18]
  reg [31:0] _RAND_117;
  reg [24:0] pages_5; // @[BTB.scala 192:18]
  reg [31:0] _RAND_118;
  reg [5:0] pageValid; // @[BTB.scala 193:22]
  reg [31:0] _RAND_119;
  reg [27:0] isValid; // @[BTB.scala 195:20]
  reg [31:0] _RAND_120;
  reg [1:0] cfiType_0; // @[BTB.scala 196:20]
  reg [31:0] _RAND_121;
  reg [1:0] cfiType_1; // @[BTB.scala 196:20]
  reg [31:0] _RAND_122;
  reg [1:0] cfiType_2; // @[BTB.scala 196:20]
  reg [31:0] _RAND_123;
  reg [1:0] cfiType_3; // @[BTB.scala 196:20]
  reg [31:0] _RAND_124;
  reg [1:0] cfiType_4; // @[BTB.scala 196:20]
  reg [31:0] _RAND_125;
  reg [1:0] cfiType_5; // @[BTB.scala 196:20]
  reg [31:0] _RAND_126;
  reg [1:0] cfiType_6; // @[BTB.scala 196:20]
  reg [31:0] _RAND_127;
  reg [1:0] cfiType_7; // @[BTB.scala 196:20]
  reg [31:0] _RAND_128;
  reg [1:0] cfiType_8; // @[BTB.scala 196:20]
  reg [31:0] _RAND_129;
  reg [1:0] cfiType_9; // @[BTB.scala 196:20]
  reg [31:0] _RAND_130;
  reg [1:0] cfiType_10; // @[BTB.scala 196:20]
  reg [31:0] _RAND_131;
  reg [1:0] cfiType_11; // @[BTB.scala 196:20]
  reg [31:0] _RAND_132;
  reg [1:0] cfiType_12; // @[BTB.scala 196:20]
  reg [31:0] _RAND_133;
  reg [1:0] cfiType_13; // @[BTB.scala 196:20]
  reg [31:0] _RAND_134;
  reg [1:0] cfiType_14; // @[BTB.scala 196:20]
  reg [31:0] _RAND_135;
  reg [1:0] cfiType_15; // @[BTB.scala 196:20]
  reg [31:0] _RAND_136;
  reg [1:0] cfiType_16; // @[BTB.scala 196:20]
  reg [31:0] _RAND_137;
  reg [1:0] cfiType_17; // @[BTB.scala 196:20]
  reg [31:0] _RAND_138;
  reg [1:0] cfiType_18; // @[BTB.scala 196:20]
  reg [31:0] _RAND_139;
  reg [1:0] cfiType_19; // @[BTB.scala 196:20]
  reg [31:0] _RAND_140;
  reg [1:0] cfiType_20; // @[BTB.scala 196:20]
  reg [31:0] _RAND_141;
  reg [1:0] cfiType_21; // @[BTB.scala 196:20]
  reg [31:0] _RAND_142;
  reg [1:0] cfiType_22; // @[BTB.scala 196:20]
  reg [31:0] _RAND_143;
  reg [1:0] cfiType_23; // @[BTB.scala 196:20]
  reg [31:0] _RAND_144;
  reg [1:0] cfiType_24; // @[BTB.scala 196:20]
  reg [31:0] _RAND_145;
  reg [1:0] cfiType_25; // @[BTB.scala 196:20]
  reg [31:0] _RAND_146;
  reg [1:0] cfiType_26; // @[BTB.scala 196:20]
  reg [31:0] _RAND_147;
  reg [1:0] cfiType_27; // @[BTB.scala 196:20]
  reg [31:0] _RAND_148;
  reg  brIdx_0; // @[BTB.scala 197:18]
  reg [31:0] _RAND_149;
  reg  brIdx_1; // @[BTB.scala 197:18]
  reg [31:0] _RAND_150;
  reg  brIdx_2; // @[BTB.scala 197:18]
  reg [31:0] _RAND_151;
  reg  brIdx_3; // @[BTB.scala 197:18]
  reg [31:0] _RAND_152;
  reg  brIdx_4; // @[BTB.scala 197:18]
  reg [31:0] _RAND_153;
  reg  brIdx_5; // @[BTB.scala 197:18]
  reg [31:0] _RAND_154;
  reg  brIdx_6; // @[BTB.scala 197:18]
  reg [31:0] _RAND_155;
  reg  brIdx_7; // @[BTB.scala 197:18]
  reg [31:0] _RAND_156;
  reg  brIdx_8; // @[BTB.scala 197:18]
  reg [31:0] _RAND_157;
  reg  brIdx_9; // @[BTB.scala 197:18]
  reg [31:0] _RAND_158;
  reg  brIdx_10; // @[BTB.scala 197:18]
  reg [31:0] _RAND_159;
  reg  brIdx_11; // @[BTB.scala 197:18]
  reg [31:0] _RAND_160;
  reg  brIdx_12; // @[BTB.scala 197:18]
  reg [31:0] _RAND_161;
  reg  brIdx_13; // @[BTB.scala 197:18]
  reg [31:0] _RAND_162;
  reg  brIdx_14; // @[BTB.scala 197:18]
  reg [31:0] _RAND_163;
  reg  brIdx_15; // @[BTB.scala 197:18]
  reg [31:0] _RAND_164;
  reg  brIdx_16; // @[BTB.scala 197:18]
  reg [31:0] _RAND_165;
  reg  brIdx_17; // @[BTB.scala 197:18]
  reg [31:0] _RAND_166;
  reg  brIdx_18; // @[BTB.scala 197:18]
  reg [31:0] _RAND_167;
  reg  brIdx_19; // @[BTB.scala 197:18]
  reg [31:0] _RAND_168;
  reg  brIdx_20; // @[BTB.scala 197:18]
  reg [31:0] _RAND_169;
  reg  brIdx_21; // @[BTB.scala 197:18]
  reg [31:0] _RAND_170;
  reg  brIdx_22; // @[BTB.scala 197:18]
  reg [31:0] _RAND_171;
  reg  brIdx_23; // @[BTB.scala 197:18]
  reg [31:0] _RAND_172;
  reg  brIdx_24; // @[BTB.scala 197:18]
  reg [31:0] _RAND_173;
  reg  brIdx_25; // @[BTB.scala 197:18]
  reg [31:0] _RAND_174;
  reg  brIdx_26; // @[BTB.scala 197:18]
  reg [31:0] _RAND_175;
  reg  brIdx_27; // @[BTB.scala 197:18]
  reg [31:0] _RAND_176;
  reg  r_btb_updatePipe_valid; // @[Valid.scala 117:22]
  reg [31:0] _RAND_177;
  reg [4:0] r_btb_updatePipe_bits_prediction_entry; // @[Reg.scala 15:16]
  reg [31:0] _RAND_178;
  reg [38:0] r_btb_updatePipe_bits_pc; // @[Reg.scala 15:16]
  reg [63:0] _RAND_179;
  reg  r_btb_updatePipe_bits_isValid; // @[Reg.scala 15:16]
  reg [31:0] _RAND_180;
  reg [38:0] r_btb_updatePipe_bits_br_pc; // @[Reg.scala 15:16]
  reg [63:0] _RAND_181;
  reg [1:0] r_btb_updatePipe_bits_cfiType; // @[Reg.scala 15:16]
  reg [31:0] _RAND_182;
  wire  _T_1; // @[BTB.scala 202:29]
  wire  _T_2; // @[BTB.scala 202:29]
  wire  _T_3; // @[BTB.scala 202:29]
  wire  _T_4; // @[BTB.scala 202:29]
  wire  _T_5; // @[BTB.scala 202:29]
  wire  _T_6; // @[BTB.scala 202:29]
  wire [5:0] _T_11; // @[Cat.scala 29:58]
  wire [5:0] pageHit; // @[BTB.scala 202:15]
  wire  _T_13; // @[BTB.scala 206:16]
  wire  _T_14; // @[BTB.scala 206:16]
  wire  _T_15; // @[BTB.scala 206:16]
  wire  _T_16; // @[BTB.scala 206:16]
  wire  _T_17; // @[BTB.scala 206:16]
  wire  _T_18; // @[BTB.scala 206:16]
  wire  _T_19; // @[BTB.scala 206:16]
  wire  _T_20; // @[BTB.scala 206:16]
  wire  _T_21; // @[BTB.scala 206:16]
  wire  _T_22; // @[BTB.scala 206:16]
  wire  _T_23; // @[BTB.scala 206:16]
  wire  _T_24; // @[BTB.scala 206:16]
  wire  _T_25; // @[BTB.scala 206:16]
  wire  _T_26; // @[BTB.scala 206:16]
  wire  _T_27; // @[BTB.scala 206:16]
  wire  _T_28; // @[BTB.scala 206:16]
  wire  _T_29; // @[BTB.scala 206:16]
  wire  _T_30; // @[BTB.scala 206:16]
  wire  _T_31; // @[BTB.scala 206:16]
  wire  _T_32; // @[BTB.scala 206:16]
  wire  _T_33; // @[BTB.scala 206:16]
  wire  _T_34; // @[BTB.scala 206:16]
  wire  _T_35; // @[BTB.scala 206:16]
  wire  _T_36; // @[BTB.scala 206:16]
  wire  _T_37; // @[BTB.scala 206:16]
  wire  _T_38; // @[BTB.scala 206:16]
  wire  _T_39; // @[BTB.scala 206:16]
  wire  _T_40; // @[BTB.scala 206:16]
  wire [6:0] _T_46; // @[Cat.scala 29:58]
  wire [13:0] _T_53; // @[Cat.scala 29:58]
  wire [6:0] _T_59; // @[Cat.scala 29:58]
  wire [27:0] _T_67; // @[Cat.scala 29:58]
  wire [27:0] idxHit; // @[BTB.scala 206:32]
  wire  _T_69; // @[BTB.scala 202:29]
  wire  _T_70; // @[BTB.scala 202:29]
  wire  _T_71; // @[BTB.scala 202:29]
  wire  _T_72; // @[BTB.scala 202:29]
  wire  _T_73; // @[BTB.scala 202:29]
  wire  _T_74; // @[BTB.scala 202:29]
  wire [5:0] _T_79; // @[Cat.scala 29:58]
  wire [5:0] updatePageHit; // @[BTB.scala 202:15]
  wire  updateHit; // @[BTB.scala 220:48]
  wire  useUpdatePageHit; // @[BTB.scala 222:40]
  wire  usePageHit; // @[BTB.scala 223:28]
  wire  doIdxPageRepl; // @[BTB.scala 224:23]
  reg [2:0] nextPageRepl; // @[BTB.scala 225:25]
  reg [31:0] _RAND_183;
  wire [5:0] _T_82; // @[Cat.scala 29:58]
  wire [7:0] _T_83; // @[OneHot.scala 58:35]
  wire [7:0] _T_84; // @[BTB.scala 226:70]
  wire [7:0] _GEN_432; // @[BTB.scala 226:65]
  wire [7:0] idxPageRepl; // @[BTB.scala 226:65]
  wire [7:0] idxPageUpdateOH; // @[BTB.scala 227:28]
  wire  _T_87; // @[OneHot.scala 32:14]
  wire [3:0] _T_88; // @[OneHot.scala 32:28]
  wire  _T_91; // @[OneHot.scala 32:14]
  wire [1:0] _T_92; // @[OneHot.scala 32:28]
  wire [2:0] idxPageUpdate; // @[Cat.scala 29:58]
  wire [7:0] idxPageReplEn; // @[BTB.scala 229:26]
  wire  samePage; // @[BTB.scala 231:45]
  wire  doTgtPageRepl; // @[BTB.scala 232:33]
  wire [5:0] _T_101; // @[Cat.scala 29:58]
  wire [7:0] tgtPageRepl; // @[BTB.scala 233:24]
  wire [7:0] _T_102; // @[BTB.scala 234:45]
  wire [7:0] _GEN_433; // @[BTB.scala 234:40]
  wire [7:0] _T_103; // @[BTB.scala 234:40]
  wire  _T_106; // @[OneHot.scala 32:14]
  wire [3:0] _T_107; // @[OneHot.scala 32:28]
  wire  _T_110; // @[OneHot.scala 32:14]
  wire [1:0] _T_111; // @[OneHot.scala 32:28]
  wire [2:0] tgtPageUpdate; // @[Cat.scala 29:58]
  wire [7:0] tgtPageReplEn; // @[BTB.scala 235:26]
  wire  _T_114; // @[BTB.scala 237:46]
  wire  _T_115; // @[BTB.scala 237:28]
  wire  _T_116; // @[BTB.scala 238:30]
  wire [1:0] _T_117; // @[BTB.scala 239:40]
  wire [2:0] _GEN_434; // @[BTB.scala 239:29]
  wire [2:0] _T_119; // @[BTB.scala 239:29]
  wire  _T_120; // @[BTB.scala 240:30]
  reg [26:0] _T_123; // @[Replacement.scala 158:30]
  reg [31:0] _RAND_184;
  wire  _T_135; // @[Replacement.scala 240:16]
  wire [1:0] _T_136; // @[Cat.scala 29:58]
  wire  _T_145; // @[Replacement.scala 240:16]
  wire [1:0] _T_146; // @[Cat.scala 29:58]
  wire  _T_152; // @[Replacement.scala 240:16]
  wire [1:0] _T_153; // @[Cat.scala 29:58]
  wire [1:0] _T_154; // @[Replacement.scala 240:16]
  wire [2:0] _T_155; // @[Cat.scala 29:58]
  wire [2:0] _T_156; // @[Replacement.scala 240:16]
  wire [3:0] _T_157; // @[Cat.scala 29:58]
  wire  _T_169; // @[Replacement.scala 240:16]
  wire [1:0] _T_170; // @[Cat.scala 29:58]
  wire  _T_176; // @[Replacement.scala 240:16]
  wire [1:0] _T_177; // @[Cat.scala 29:58]
  wire [1:0] _T_178; // @[Replacement.scala 240:16]
  wire [2:0] _T_179; // @[Cat.scala 29:58]
  wire  _T_188; // @[Replacement.scala 240:16]
  wire [1:0] _T_189; // @[Cat.scala 29:58]
  wire  _T_195; // @[Replacement.scala 240:16]
  wire [1:0] _T_196; // @[Cat.scala 29:58]
  wire [1:0] _T_197; // @[Replacement.scala 240:16]
  wire [2:0] _T_198; // @[Cat.scala 29:58]
  wire [2:0] _T_199; // @[Replacement.scala 240:16]
  wire [3:0] _T_200; // @[Cat.scala 29:58]
  wire [3:0] _T_201; // @[Replacement.scala 240:16]
  wire [4:0] _T_202; // @[Cat.scala 29:58]
  wire [4:0] waddr; // @[BTB.scala 244:18]
  reg  r_respPipe_valid; // @[Valid.scala 117:22]
  reg [31:0] _RAND_185;
  reg  r_respPipe_bits_taken; // @[Reg.scala 15:16]
  reg [31:0] _RAND_186;
  reg [4:0] r_respPipe_bits_entry; // @[Reg.scala 15:16]
  reg [31:0] _RAND_187;
  wire  _T_203; // @[BTB.scala 246:22]
  wire  _T_204; // @[BTB.scala 246:43]
  wire [4:0] _T_205; // @[BTB.scala 247:20]
  wire  _T_224; // @[Replacement.scala 193:16]
  wire  _T_228; // @[Replacement.scala 196:16]
  wire [2:0] _T_230; // @[Cat.scala 29:58]
  wire [2:0] _T_231; // @[Replacement.scala 193:16]
  wire  _T_245; // @[Replacement.scala 193:16]
  wire  _T_249; // @[Replacement.scala 196:16]
  wire [2:0] _T_251; // @[Cat.scala 29:58]
  wire [2:0] _T_252; // @[Replacement.scala 193:16]
  wire  _T_261; // @[Replacement.scala 193:16]
  wire  _T_265; // @[Replacement.scala 196:16]
  wire [2:0] _T_267; // @[Cat.scala 29:58]
  wire [2:0] _T_268; // @[Replacement.scala 196:16]
  wire [6:0] _T_270; // @[Cat.scala 29:58]
  wire [6:0] _T_271; // @[Replacement.scala 196:16]
  wire [10:0] _T_273; // @[Cat.scala 29:58]
  wire [10:0] _T_274; // @[Replacement.scala 193:16]
  wire  _T_293; // @[Replacement.scala 193:16]
  wire  _T_297; // @[Replacement.scala 196:16]
  wire [2:0] _T_299; // @[Cat.scala 29:58]
  wire [2:0] _T_300; // @[Replacement.scala 193:16]
  wire  _T_309; // @[Replacement.scala 193:16]
  wire  _T_313; // @[Replacement.scala 196:16]
  wire [2:0] _T_315; // @[Cat.scala 29:58]
  wire [2:0] _T_316; // @[Replacement.scala 196:16]
  wire [6:0] _T_318; // @[Cat.scala 29:58]
  wire [6:0] _T_319; // @[Replacement.scala 193:16]
  wire  _T_333; // @[Replacement.scala 193:16]
  wire  _T_337; // @[Replacement.scala 196:16]
  wire [2:0] _T_339; // @[Cat.scala 29:58]
  wire [2:0] _T_340; // @[Replacement.scala 193:16]
  wire  _T_349; // @[Replacement.scala 193:16]
  wire  _T_353; // @[Replacement.scala 196:16]
  wire [2:0] _T_355; // @[Cat.scala 29:58]
  wire [2:0] _T_356; // @[Replacement.scala 196:16]
  wire [6:0] _T_358; // @[Cat.scala 29:58]
  wire [6:0] _T_359; // @[Replacement.scala 196:16]
  wire [14:0] _T_361; // @[Cat.scala 29:58]
  wire [14:0] _T_362; // @[Replacement.scala 196:16]
  wire [26:0] _T_364; // @[Cat.scala 29:58]
  wire [31:0] _T_365; // @[OneHot.scala 58:35]
  wire [3:0] _T_368; // @[BTB.scala 254:38]
  wire [31:0] _GEN_435; // @[BTB.scala 257:55]
  wire [31:0] _T_369; // @[BTB.scala 257:55]
  wire [31:0] _T_371; // @[BTB.scala 257:71]
  wire [31:0] _T_372; // @[BTB.scala 257:19]
  wire [7:0] _T_376; // @[BTB.scala 268:24]
  wire [7:0] _T_383; // @[BTB.scala 270:24]
  wire [7:0] _GEN_437; // @[BTB.scala 272:28]
  wire [7:0] _T_390; // @[BTB.scala 272:28]
  wire [7:0] _T_391; // @[BTB.scala 272:44]
  wire [31:0] _GEN_338; // @[BTB.scala 250:29]
  wire [7:0] _GEN_373; // @[BTB.scala 250:29]
  wire [6:0] _T_392; // @[BTB.scala 275:29]
  wire [2:0] _T_421; // @[Mux.scala 27:72]
  wire [2:0] _T_422; // @[Mux.scala 27:72]
  wire [2:0] _T_423; // @[Mux.scala 27:72]
  wire [2:0] _T_424; // @[Mux.scala 27:72]
  wire [2:0] _T_425; // @[Mux.scala 27:72]
  wire [2:0] _T_426; // @[Mux.scala 27:72]
  wire [2:0] _T_427; // @[Mux.scala 27:72]
  wire [2:0] _T_428; // @[Mux.scala 27:72]
  wire [2:0] _T_429; // @[Mux.scala 27:72]
  wire [2:0] _T_430; // @[Mux.scala 27:72]
  wire [2:0] _T_431; // @[Mux.scala 27:72]
  wire [2:0] _T_432; // @[Mux.scala 27:72]
  wire [2:0] _T_433; // @[Mux.scala 27:72]
  wire [2:0] _T_434; // @[Mux.scala 27:72]
  wire [2:0] _T_435; // @[Mux.scala 27:72]
  wire [2:0] _T_436; // @[Mux.scala 27:72]
  wire [2:0] _T_437; // @[Mux.scala 27:72]
  wire [2:0] _T_438; // @[Mux.scala 27:72]
  wire [2:0] _T_439; // @[Mux.scala 27:72]
  wire [2:0] _T_440; // @[Mux.scala 27:72]
  wire [2:0] _T_441; // @[Mux.scala 27:72]
  wire [2:0] _T_442; // @[Mux.scala 27:72]
  wire [2:0] _T_443; // @[Mux.scala 27:72]
  wire [2:0] _T_444; // @[Mux.scala 27:72]
  wire [2:0] _T_445; // @[Mux.scala 27:72]
  wire [2:0] _T_446; // @[Mux.scala 27:72]
  wire [2:0] _T_447; // @[Mux.scala 27:72]
  wire [2:0] _T_448; // @[Mux.scala 27:72]
  wire [2:0] _T_449; // @[Mux.scala 27:72]
  wire [2:0] _T_450; // @[Mux.scala 27:72]
  wire [2:0] _T_451; // @[Mux.scala 27:72]
  wire [2:0] _T_452; // @[Mux.scala 27:72]
  wire [2:0] _T_453; // @[Mux.scala 27:72]
  wire [2:0] _T_454; // @[Mux.scala 27:72]
  wire [2:0] _T_455; // @[Mux.scala 27:72]
  wire [2:0] _T_456; // @[Mux.scala 27:72]
  wire [2:0] _T_457; // @[Mux.scala 27:72]
  wire [2:0] _T_458; // @[Mux.scala 27:72]
  wire [2:0] _T_459; // @[Mux.scala 27:72]
  wire [2:0] _T_460; // @[Mux.scala 27:72]
  wire [2:0] _T_461; // @[Mux.scala 27:72]
  wire [2:0] _T_462; // @[Mux.scala 27:72]
  wire [2:0] _T_463; // @[Mux.scala 27:72]
  wire [2:0] _T_464; // @[Mux.scala 27:72]
  wire [2:0] _T_465; // @[Mux.scala 27:72]
  wire [2:0] _T_466; // @[Mux.scala 27:72]
  wire [2:0] _T_467; // @[Mux.scala 27:72]
  wire [2:0] _T_468; // @[Mux.scala 27:72]
  wire [2:0] _T_469; // @[Mux.scala 27:72]
  wire [2:0] _T_470; // @[Mux.scala 27:72]
  wire [2:0] _T_471; // @[Mux.scala 27:72]
  wire [2:0] _T_472; // @[Mux.scala 27:72]
  wire [2:0] _T_473; // @[Mux.scala 27:72]
  wire [2:0] _T_474; // @[Mux.scala 27:72]
  wire [2:0] _T_475; // @[Mux.scala 27:72]
  wire [6:0] _T_477; // @[BTB.scala 275:34]
  wire [2:0] _T_507; // @[Mux.scala 27:72]
  wire [2:0] _T_508; // @[Mux.scala 27:72]
  wire [2:0] _T_509; // @[Mux.scala 27:72]
  wire [2:0] _T_510; // @[Mux.scala 27:72]
  wire [2:0] _T_511; // @[Mux.scala 27:72]
  wire [2:0] _T_512; // @[Mux.scala 27:72]
  wire [2:0] _T_513; // @[Mux.scala 27:72]
  wire [2:0] _T_514; // @[Mux.scala 27:72]
  wire [2:0] _T_515; // @[Mux.scala 27:72]
  wire [2:0] _T_516; // @[Mux.scala 27:72]
  wire [2:0] _T_517; // @[Mux.scala 27:72]
  wire [2:0] _T_518; // @[Mux.scala 27:72]
  wire [2:0] _T_519; // @[Mux.scala 27:72]
  wire [2:0] _T_520; // @[Mux.scala 27:72]
  wire [2:0] _T_521; // @[Mux.scala 27:72]
  wire [2:0] _T_522; // @[Mux.scala 27:72]
  wire [2:0] _T_523; // @[Mux.scala 27:72]
  wire [2:0] _T_524; // @[Mux.scala 27:72]
  wire [2:0] _T_525; // @[Mux.scala 27:72]
  wire [2:0] _T_526; // @[Mux.scala 27:72]
  wire [2:0] _T_527; // @[Mux.scala 27:72]
  wire [2:0] _T_528; // @[Mux.scala 27:72]
  wire [2:0] _T_529; // @[Mux.scala 27:72]
  wire [2:0] _T_530; // @[Mux.scala 27:72]
  wire [2:0] _T_531; // @[Mux.scala 27:72]
  wire [2:0] _T_532; // @[Mux.scala 27:72]
  wire [2:0] _T_533; // @[Mux.scala 27:72]
  wire [2:0] _T_534; // @[Mux.scala 27:72]
  wire [2:0] _T_535; // @[Mux.scala 27:72]
  wire [2:0] _T_536; // @[Mux.scala 27:72]
  wire [2:0] _T_537; // @[Mux.scala 27:72]
  wire [2:0] _T_538; // @[Mux.scala 27:72]
  wire [2:0] _T_539; // @[Mux.scala 27:72]
  wire [2:0] _T_540; // @[Mux.scala 27:72]
  wire [2:0] _T_541; // @[Mux.scala 27:72]
  wire [2:0] _T_542; // @[Mux.scala 27:72]
  wire [2:0] _T_543; // @[Mux.scala 27:72]
  wire [2:0] _T_544; // @[Mux.scala 27:72]
  wire [2:0] _T_545; // @[Mux.scala 27:72]
  wire [2:0] _T_546; // @[Mux.scala 27:72]
  wire [2:0] _T_547; // @[Mux.scala 27:72]
  wire [2:0] _T_548; // @[Mux.scala 27:72]
  wire [2:0] _T_549; // @[Mux.scala 27:72]
  wire [2:0] _T_550; // @[Mux.scala 27:72]
  wire [2:0] _T_551; // @[Mux.scala 27:72]
  wire [2:0] _T_552; // @[Mux.scala 27:72]
  wire [2:0] _T_553; // @[Mux.scala 27:72]
  wire [2:0] _T_554; // @[Mux.scala 27:72]
  wire [2:0] _T_555; // @[Mux.scala 27:72]
  wire [2:0] _T_556; // @[Mux.scala 27:72]
  wire [2:0] _T_557; // @[Mux.scala 27:72]
  wire [2:0] _T_558; // @[Mux.scala 27:72]
  wire [2:0] _T_559; // @[Mux.scala 27:72]
  wire [2:0] _T_560; // @[Mux.scala 27:72]
  wire [2:0] _T_561; // @[Mux.scala 27:72]
  wire [12:0] _T_591; // @[Mux.scala 27:72]
  wire [12:0] _T_592; // @[Mux.scala 27:72]
  wire [12:0] _T_593; // @[Mux.scala 27:72]
  wire [12:0] _T_594; // @[Mux.scala 27:72]
  wire [12:0] _T_595; // @[Mux.scala 27:72]
  wire [12:0] _T_596; // @[Mux.scala 27:72]
  wire [12:0] _T_597; // @[Mux.scala 27:72]
  wire [12:0] _T_598; // @[Mux.scala 27:72]
  wire [12:0] _T_599; // @[Mux.scala 27:72]
  wire [12:0] _T_600; // @[Mux.scala 27:72]
  wire [12:0] _T_601; // @[Mux.scala 27:72]
  wire [12:0] _T_602; // @[Mux.scala 27:72]
  wire [12:0] _T_603; // @[Mux.scala 27:72]
  wire [12:0] _T_604; // @[Mux.scala 27:72]
  wire [12:0] _T_605; // @[Mux.scala 27:72]
  wire [12:0] _T_606; // @[Mux.scala 27:72]
  wire [12:0] _T_607; // @[Mux.scala 27:72]
  wire [12:0] _T_608; // @[Mux.scala 27:72]
  wire [12:0] _T_609; // @[Mux.scala 27:72]
  wire [12:0] _T_610; // @[Mux.scala 27:72]
  wire [12:0] _T_611; // @[Mux.scala 27:72]
  wire [12:0] _T_612; // @[Mux.scala 27:72]
  wire [12:0] _T_613; // @[Mux.scala 27:72]
  wire [12:0] _T_614; // @[Mux.scala 27:72]
  wire [12:0] _T_615; // @[Mux.scala 27:72]
  wire [12:0] _T_616; // @[Mux.scala 27:72]
  wire [12:0] _T_617; // @[Mux.scala 27:72]
  wire [12:0] _T_618; // @[Mux.scala 27:72]
  wire [12:0] _T_619; // @[Mux.scala 27:72]
  wire [12:0] _T_620; // @[Mux.scala 27:72]
  wire [12:0] _T_621; // @[Mux.scala 27:72]
  wire [12:0] _T_622; // @[Mux.scala 27:72]
  wire [12:0] _T_623; // @[Mux.scala 27:72]
  wire [12:0] _T_624; // @[Mux.scala 27:72]
  wire [12:0] _T_625; // @[Mux.scala 27:72]
  wire [12:0] _T_626; // @[Mux.scala 27:72]
  wire [12:0] _T_627; // @[Mux.scala 27:72]
  wire [12:0] _T_628; // @[Mux.scala 27:72]
  wire [12:0] _T_629; // @[Mux.scala 27:72]
  wire [12:0] _T_630; // @[Mux.scala 27:72]
  wire [12:0] _T_631; // @[Mux.scala 27:72]
  wire [12:0] _T_632; // @[Mux.scala 27:72]
  wire [12:0] _T_633; // @[Mux.scala 27:72]
  wire [12:0] _T_634; // @[Mux.scala 27:72]
  wire [12:0] _T_635; // @[Mux.scala 27:72]
  wire [12:0] _T_636; // @[Mux.scala 27:72]
  wire [12:0] _T_637; // @[Mux.scala 27:72]
  wire [12:0] _T_638; // @[Mux.scala 27:72]
  wire [12:0] _T_639; // @[Mux.scala 27:72]
  wire [12:0] _T_640; // @[Mux.scala 27:72]
  wire [12:0] _T_641; // @[Mux.scala 27:72]
  wire [12:0] _T_642; // @[Mux.scala 27:72]
  wire [12:0] _T_643; // @[Mux.scala 27:72]
  wire [12:0] _T_644; // @[Mux.scala 27:72]
  wire [12:0] _T_645; // @[Mux.scala 27:72]
  wire [13:0] _T_647; // @[BTB.scala 277:82]
  wire [24:0] _GEN_375; // @[Cat.scala 29:58]
  wire [24:0] _GEN_376; // @[Cat.scala 29:58]
  wire [24:0] _GEN_377; // @[Cat.scala 29:58]
  wire [24:0] _GEN_378; // @[Cat.scala 29:58]
  wire [24:0] _GEN_379; // @[Cat.scala 29:58]
  wire [38:0] _T_648; // @[Cat.scala 29:58]
  wire  _T_651; // @[OneHot.scala 32:14]
  wire [15:0] _GEN_438; // @[OneHot.scala 32:28]
  wire [15:0] _T_652; // @[OneHot.scala 32:28]
  wire  _T_655; // @[OneHot.scala 32:14]
  wire [7:0] _T_656; // @[OneHot.scala 32:28]
  wire  _T_659; // @[OneHot.scala 32:14]
  wire [3:0] _T_660; // @[OneHot.scala 32:28]
  wire  _T_663; // @[OneHot.scala 32:14]
  wire [1:0] _T_664; // @[OneHot.scala 32:28]
  wire [3:0] _T_668; // @[Cat.scala 29:58]
  wire  _T_698; // @[Mux.scala 27:72]
  wire  _T_699; // @[Mux.scala 27:72]
  wire  _T_700; // @[Mux.scala 27:72]
  wire  _T_701; // @[Mux.scala 27:72]
  wire  _T_702; // @[Mux.scala 27:72]
  wire  _T_703; // @[Mux.scala 27:72]
  wire  _T_704; // @[Mux.scala 27:72]
  wire  _T_705; // @[Mux.scala 27:72]
  wire  _T_706; // @[Mux.scala 27:72]
  wire  _T_707; // @[Mux.scala 27:72]
  wire  _T_708; // @[Mux.scala 27:72]
  wire  _T_709; // @[Mux.scala 27:72]
  wire  _T_710; // @[Mux.scala 27:72]
  wire  _T_711; // @[Mux.scala 27:72]
  wire  _T_712; // @[Mux.scala 27:72]
  wire  _T_713; // @[Mux.scala 27:72]
  wire  _T_714; // @[Mux.scala 27:72]
  wire  _T_715; // @[Mux.scala 27:72]
  wire  _T_716; // @[Mux.scala 27:72]
  wire  _T_717; // @[Mux.scala 27:72]
  wire  _T_718; // @[Mux.scala 27:72]
  wire  _T_719; // @[Mux.scala 27:72]
  wire  _T_720; // @[Mux.scala 27:72]
  wire  _T_721; // @[Mux.scala 27:72]
  wire  _T_722; // @[Mux.scala 27:72]
  wire  _T_723; // @[Mux.scala 27:72]
  wire  _T_724; // @[Mux.scala 27:72]
  wire  _T_725; // @[Mux.scala 27:72]
  wire  _T_726; // @[Mux.scala 27:72]
  wire  _T_727; // @[Mux.scala 27:72]
  wire  _T_728; // @[Mux.scala 27:72]
  wire  _T_729; // @[Mux.scala 27:72]
  wire  _T_730; // @[Mux.scala 27:72]
  wire  _T_731; // @[Mux.scala 27:72]
  wire  _T_732; // @[Mux.scala 27:72]
  wire  _T_733; // @[Mux.scala 27:72]
  wire  _T_734; // @[Mux.scala 27:72]
  wire  _T_735; // @[Mux.scala 27:72]
  wire  _T_736; // @[Mux.scala 27:72]
  wire  _T_737; // @[Mux.scala 27:72]
  wire  _T_738; // @[Mux.scala 27:72]
  wire  _T_739; // @[Mux.scala 27:72]
  wire  _T_740; // @[Mux.scala 27:72]
  wire  _T_741; // @[Mux.scala 27:72]
  wire  _T_742; // @[Mux.scala 27:72]
  wire  _T_743; // @[Mux.scala 27:72]
  wire  _T_744; // @[Mux.scala 27:72]
  wire  _T_745; // @[Mux.scala 27:72]
  wire  _T_746; // @[Mux.scala 27:72]
  wire  _T_747; // @[Mux.scala 27:72]
  wire  _T_748; // @[Mux.scala 27:72]
  wire  _T_749; // @[Mux.scala 27:72]
  wire  _T_750; // @[Mux.scala 27:72]
  wire  _T_751; // @[Mux.scala 27:72]
  wire  _T_855; // @[Misc.scala 182:16]
  wire  _T_857; // @[Misc.scala 182:61]
  wire  _T_859; // @[Misc.scala 182:16]
  wire  _T_861; // @[Misc.scala 182:61]
  wire  _T_862; // @[Misc.scala 182:49]
  wire  _T_869; // @[Misc.scala 182:16]
  wire  _T_871; // @[Misc.scala 182:61]
  wire  _T_878; // @[Misc.scala 182:16]
  wire  _T_880; // @[Misc.scala 182:61]
  wire  _T_882; // @[Misc.scala 182:16]
  wire  _T_883; // @[Misc.scala 182:37]
  wire  _T_884; // @[Misc.scala 182:61]
  wire  _T_885; // @[Misc.scala 182:49]
  wire  _T_886; // @[Misc.scala 182:16]
  wire  _T_887; // @[Misc.scala 182:37]
  wire  _T_888; // @[Misc.scala 182:61]
  wire  _T_889; // @[Misc.scala 182:49]
  wire  _T_899; // @[Misc.scala 182:16]
  wire  _T_901; // @[Misc.scala 182:61]
  wire  _T_903; // @[Misc.scala 182:16]
  wire  _T_905; // @[Misc.scala 182:61]
  wire  _T_906; // @[Misc.scala 182:49]
  wire  _T_913; // @[Misc.scala 182:16]
  wire  _T_915; // @[Misc.scala 182:61]
  wire  _T_922; // @[Misc.scala 182:16]
  wire  _T_924; // @[Misc.scala 182:61]
  wire  _T_926; // @[Misc.scala 182:16]
  wire  _T_927; // @[Misc.scala 182:37]
  wire  _T_928; // @[Misc.scala 182:61]
  wire  _T_929; // @[Misc.scala 182:49]
  wire  _T_930; // @[Misc.scala 182:16]
  wire  _T_931; // @[Misc.scala 182:37]
  wire  _T_932; // @[Misc.scala 182:61]
  wire  _T_933; // @[Misc.scala 182:49]
  wire  _T_934; // @[Misc.scala 182:16]
  wire  _T_935; // @[Misc.scala 182:37]
  wire  _T_936; // @[Misc.scala 182:61]
  wire  _T_937; // @[Misc.scala 182:49]
  wire  _T_948; // @[Misc.scala 182:16]
  wire  _T_950; // @[Misc.scala 182:61]
  wire  _T_952; // @[Misc.scala 182:16]
  wire  _T_954; // @[Misc.scala 182:61]
  wire  _T_955; // @[Misc.scala 182:49]
  wire  _T_962; // @[Misc.scala 182:16]
  wire  _T_964; // @[Misc.scala 182:61]
  wire  _T_971; // @[Misc.scala 182:16]
  wire  _T_973; // @[Misc.scala 182:61]
  wire  _T_975; // @[Misc.scala 182:16]
  wire  _T_976; // @[Misc.scala 182:37]
  wire  _T_977; // @[Misc.scala 182:61]
  wire  _T_978; // @[Misc.scala 182:49]
  wire  _T_979; // @[Misc.scala 182:16]
  wire  _T_980; // @[Misc.scala 182:37]
  wire  _T_981; // @[Misc.scala 182:61]
  wire  _T_982; // @[Misc.scala 182:49]
  wire  _T_992; // @[Misc.scala 182:16]
  wire  _T_994; // @[Misc.scala 182:61]
  wire  _T_996; // @[Misc.scala 182:16]
  wire  _T_998; // @[Misc.scala 182:61]
  wire  _T_999; // @[Misc.scala 182:49]
  wire  _T_1006; // @[Misc.scala 182:16]
  wire  _T_1008; // @[Misc.scala 182:61]
  wire  _T_1015; // @[Misc.scala 182:16]
  wire  _T_1017; // @[Misc.scala 182:61]
  wire  _T_1019; // @[Misc.scala 182:16]
  wire  _T_1020; // @[Misc.scala 182:37]
  wire  _T_1021; // @[Misc.scala 182:61]
  wire  _T_1022; // @[Misc.scala 182:49]
  wire  _T_1023; // @[Misc.scala 182:16]
  wire  _T_1024; // @[Misc.scala 182:37]
  wire  _T_1025; // @[Misc.scala 182:61]
  wire  _T_1026; // @[Misc.scala 182:49]
  wire  _T_1027; // @[Misc.scala 182:16]
  wire  _T_1028; // @[Misc.scala 182:37]
  wire  _T_1029; // @[Misc.scala 182:61]
  wire  _T_1030; // @[Misc.scala 182:49]
  wire  _T_1032; // @[Misc.scala 182:37]
  wire  _T_1033; // @[Misc.scala 182:61]
  wire  _T_1034; // @[Misc.scala 182:49]
  wire [27:0] _T_1036; // @[BTB.scala 285:24]
  wire [31:0] _GEN_380; // @[BTB.scala 284:37]
  wire [31:0] _GEN_381; // @[BTB.scala 287:19]
  reg [7:0] _T_1038; // @[BTB.scala 114:20]
  reg [31:0] _RAND_188;
  wire  _T_1039; // @[BTB.scala 293:44]
  wire  _T_1040; // @[BTB.scala 293:44]
  wire  _T_1041; // @[BTB.scala 293:44]
  wire  _T_1042; // @[BTB.scala 293:44]
  wire  _T_1043; // @[BTB.scala 293:44]
  wire  _T_1044; // @[BTB.scala 293:44]
  wire  _T_1045; // @[BTB.scala 293:44]
  wire  _T_1046; // @[BTB.scala 293:44]
  wire  _T_1047; // @[BTB.scala 293:44]
  wire  _T_1048; // @[BTB.scala 293:44]
  wire  _T_1049; // @[BTB.scala 293:44]
  wire  _T_1050; // @[BTB.scala 293:44]
  wire  _T_1051; // @[BTB.scala 293:44]
  wire  _T_1052; // @[BTB.scala 293:44]
  wire  _T_1053; // @[BTB.scala 293:44]
  wire  _T_1054; // @[BTB.scala 293:44]
  wire  _T_1055; // @[BTB.scala 293:44]
  wire  _T_1056; // @[BTB.scala 293:44]
  wire  _T_1057; // @[BTB.scala 293:44]
  wire  _T_1058; // @[BTB.scala 293:44]
  wire  _T_1059; // @[BTB.scala 293:44]
  wire  _T_1060; // @[BTB.scala 293:44]
  wire  _T_1061; // @[BTB.scala 293:44]
  wire  _T_1062; // @[BTB.scala 293:44]
  wire  _T_1063; // @[BTB.scala 293:44]
  wire  _T_1064; // @[BTB.scala 293:44]
  wire  _T_1065; // @[BTB.scala 293:44]
  wire  _T_1066; // @[BTB.scala 293:44]
  wire [6:0] _T_1072; // @[Cat.scala 29:58]
  wire [13:0] _T_1079; // @[Cat.scala 29:58]
  wire [6:0] _T_1085; // @[Cat.scala 29:58]
  wire [27:0] _T_1093; // @[Cat.scala 29:58]
  wire [27:0] _T_1094; // @[BTB.scala 293:28]
  wire  _T_1095; // @[BTB.scala 293:72]
  wire [8:0] _GEN_439; // @[BTB.scala 87:42]
  wire [8:0] _T_1101; // @[BTB.scala 87:42]
  wire [15:0] _T_1102; // @[BTB.scala 83:12]
  wire [8:0] _T_1104; // @[BTB.scala 89:44]
  wire [7:0] _T_1109; // @[Cat.scala 29:58]
  wire [8:0] _GEN_440; // @[BTB.scala 87:42]
  wire [8:0] _T_1114; // @[BTB.scala 87:42]
  wire [15:0] _T_1115; // @[BTB.scala 83:12]
  wire [8:0] _T_1117; // @[BTB.scala 89:44]
  wire [7:0] _T_1121; // @[Cat.scala 29:58]
  wire  _T_1096_value; // @[BTB.scala 92:19 BTB.scala 93:15]
  wire  _T_1124; // @[BTB.scala 308:22]
  reg [2:0] _T_1125; // @[BTB.scala 57:26]
  reg [31:0] _RAND_189;
  reg [2:0] _T_1126; // @[BTB.scala 58:24]
  reg [31:0] _RAND_190;
  reg [38:0] _T_1127_0; // @[BTB.scala 59:26]
  reg [63:0] _RAND_191;
  reg [38:0] _T_1127_1; // @[BTB.scala 59:26]
  reg [63:0] _RAND_192;
  reg [38:0] _T_1127_2; // @[BTB.scala 59:26]
  reg [63:0] _RAND_193;
  reg [38:0] _T_1127_3; // @[BTB.scala 59:26]
  reg [63:0] _RAND_194;
  reg [38:0] _T_1127_4; // @[BTB.scala 59:26]
  reg [63:0] _RAND_195;
  reg [38:0] _T_1127_5; // @[BTB.scala 59:26]
  reg [63:0] _RAND_196;
  wire  _T_1128; // @[BTB.scala 314:42]
  wire  _T_1129; // @[BTB.scala 314:42]
  wire  _T_1130; // @[BTB.scala 314:42]
  wire  _T_1131; // @[BTB.scala 314:42]
  wire  _T_1132; // @[BTB.scala 314:42]
  wire  _T_1133; // @[BTB.scala 314:42]
  wire  _T_1134; // @[BTB.scala 314:42]
  wire  _T_1135; // @[BTB.scala 314:42]
  wire  _T_1136; // @[BTB.scala 314:42]
  wire  _T_1137; // @[BTB.scala 314:42]
  wire  _T_1138; // @[BTB.scala 314:42]
  wire  _T_1139; // @[BTB.scala 314:42]
  wire  _T_1140; // @[BTB.scala 314:42]
  wire  _T_1141; // @[BTB.scala 314:42]
  wire  _T_1142; // @[BTB.scala 314:42]
  wire  _T_1143; // @[BTB.scala 314:42]
  wire  _T_1144; // @[BTB.scala 314:42]
  wire  _T_1145; // @[BTB.scala 314:42]
  wire  _T_1146; // @[BTB.scala 314:42]
  wire  _T_1147; // @[BTB.scala 314:42]
  wire  _T_1148; // @[BTB.scala 314:42]
  wire  _T_1149; // @[BTB.scala 314:42]
  wire  _T_1150; // @[BTB.scala 314:42]
  wire  _T_1151; // @[BTB.scala 314:42]
  wire  _T_1152; // @[BTB.scala 314:42]
  wire  _T_1153; // @[BTB.scala 314:42]
  wire  _T_1154; // @[BTB.scala 314:42]
  wire  _T_1155; // @[BTB.scala 314:42]
  wire [6:0] _T_1161; // @[Cat.scala 29:58]
  wire [13:0] _T_1168; // @[Cat.scala 29:58]
  wire [6:0] _T_1174; // @[Cat.scala 29:58]
  wire [27:0] _T_1182; // @[Cat.scala 29:58]
  wire [27:0] _T_1183; // @[BTB.scala 314:26]
  wire  _T_1184; // @[BTB.scala 314:67]
  wire  _T_1185; // @[BTB.scala 55:29]
  wire [38:0] _GEN_399; // @[BTB.scala 316:22]
  wire [38:0] _GEN_400; // @[BTB.scala 316:22]
  wire [38:0] _GEN_401; // @[BTB.scala 316:22]
  wire [38:0] _GEN_402; // @[BTB.scala 316:22]
  wire [38:0] _GEN_403; // @[BTB.scala 316:22]
  wire  _T_1189; // @[BTB.scala 317:24]
  wire  _T_1190; // @[BTB.scala 321:40]
  wire  _T_1191; // @[BTB.scala 44:17]
  wire [2:0] _T_1193; // @[BTB.scala 44:42]
  wire  _T_1194; // @[BTB.scala 45:49]
  wire [2:0] _T_1197; // @[BTB.scala 45:62]
  wire [2:0] _T_1198; // @[BTB.scala 45:22]
  wire  _T_1199; // @[BTB.scala 323:46]
  wire [2:0] _T_1203; // @[BTB.scala 51:20]
  wire  _T_1204; // @[BTB.scala 52:42]
  wire [2:0] _T_1207; // @[BTB.scala 52:50]
  reg [19:0] BTB_state; // @[Register tracking BTB state]
  reg [31:0] _RAND_197;
  reg  BTB_cov [0:1048575]; // @[Coverage map for BTB]
  reg [31:0] _RAND_198;
  wire  BTB_cov_read_data; // @[Coverage map for BTB]
  wire [19:0] BTB_cov_read_addr; // @[Coverage map for BTB]
  wire  BTB_cov_write_data; // @[Coverage map for BTB]
  wire [19:0] BTB_cov_write_addr; // @[Coverage map for BTB]
  wire  BTB_cov_write_mask; // @[Coverage map for BTB]
  wire  BTB_cov_write_en; // @[Coverage map for BTB]
  reg [29:0] BTB_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_199;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire  mux_cond_6;
  wire  mux_cond_7;
  wire  mux_cond_8;
  wire  mux_cond_9;
  wire  mux_cond_10;
  wire  mux_cond_11;
  wire  mux_cond_12;
  wire  mux_cond_13;
  wire  mux_cond_14;
  wire  mux_cond_15;
  wire  mux_cond_16;
  wire  mux_cond_17;
  wire  mux_cond_18;
  wire  mux_cond_19;
  wire  mux_cond_20;
  wire  mux_cond_21;
  wire  mux_cond_22;
  wire  mux_cond_23;
  wire  mux_cond_24;
  wire  mux_cond_25;
  wire  mux_cond_26;
  wire  mux_cond_27;
  wire  mux_cond_28;
  wire [6:0] r_respPipe_bits_taken_shl;
  wire [19:0] r_respPipe_bits_taken_pad;
  wire [16:0] r_btb_updatePipe_valid_shl;
  wire [19:0] r_btb_updatePipe_valid_pad;
  wire [14:0] r_respPipe_valid_shl;
  wire [19:0] r_respPipe_valid_pad;
  wire [17:0] pageValid_shl;
  wire [19:0] pageValid_pad;
  wire [17:0] _T_1125_shl;
  wire [19:0] _T_1125_pad;
  wire [10:0] r_btb_updatePipe_bits_isValid_shl;
  wire [19:0] r_btb_updatePipe_bits_isValid_pad;
  wire [14:0] nextPageRepl_shl;
  wire [19:0] nextPageRepl_pad;
  wire [18:0] _T_1126_shl;
  wire [19:0] _T_1126_pad;
  wire [17:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [2:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [3:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [5:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [13:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [18:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [9:0] mux_cond_6_shl;
  wire [19:0] mux_cond_6_pad;
  wire [8:0] mux_cond_7_shl;
  wire [19:0] mux_cond_7_pad;
  wire [12:0] mux_cond_8_shl;
  wire [19:0] mux_cond_8_pad;
  wire [8:0] mux_cond_9_shl;
  wire [19:0] mux_cond_9_pad;
  wire [13:0] mux_cond_10_shl;
  wire [19:0] mux_cond_10_pad;
  wire [18:0] mux_cond_11_shl;
  wire [19:0] mux_cond_11_pad;
  wire [17:0] mux_cond_12_shl;
  wire [19:0] mux_cond_12_pad;
  wire [16:0] mux_cond_13_shl;
  wire [19:0] mux_cond_13_pad;
  wire [15:0] mux_cond_14_shl;
  wire [19:0] mux_cond_14_pad;
  wire [1:0] mux_cond_15_shl;
  wire [19:0] mux_cond_15_pad;
  wire [5:0] mux_cond_16_shl;
  wire [19:0] mux_cond_16_pad;
  wire [3:0] mux_cond_17_shl;
  wire [19:0] mux_cond_17_pad;
  wire [9:0] mux_cond_18_shl;
  wire [19:0] mux_cond_18_pad;
  wire [7:0] mux_cond_19_shl;
  wire [19:0] mux_cond_19_pad;
  wire [18:0] mux_cond_20_shl;
  wire [19:0] mux_cond_20_pad;
  wire [4:0] mux_cond_21_shl;
  wire [19:0] mux_cond_21_pad;
  wire [16:0] mux_cond_22_shl;
  wire [19:0] mux_cond_22_pad;
  wire  mux_cond_23_shl;
  wire [19:0] mux_cond_23_pad;
  wire [19:0] mux_cond_24_shl;
  wire [19:0] mux_cond_24_pad;
  wire [5:0] mux_cond_25_shl;
  wire [19:0] mux_cond_25_pad;
  wire [15:0] mux_cond_26_shl;
  wire [19:0] mux_cond_26_pad;
  wire [9:0] mux_cond_27_shl;
  wire [19:0] mux_cond_27_pad;
  wire [12:0] mux_cond_28_shl;
  wire [19:0] mux_cond_28_pad;
  wire [13:0] cfiType_4_shl;
  wire [19:0] cfiType_4_pad;
  wire [9:0] tgtPages_20_shl;
  wire [19:0] tgtPages_20_pad;
  wire [9:0] tgtPages_17_shl;
  wire [19:0] tgtPages_17_pad;
  wire [9:0] tgtPages_3_shl;
  wire [19:0] tgtPages_3_pad;
  wire [13:0] cfiType_1_shl;
  wire [19:0] cfiType_1_pad;
  wire [9:0] tgtPages_2_shl;
  wire [19:0] tgtPages_2_pad;
  wire [13:0] cfiType_18_shl;
  wire [19:0] cfiType_18_pad;
  wire [9:0] tgtPages_26_shl;
  wire [19:0] tgtPages_26_pad;
  wire [13:0] cfiType_20_shl;
  wire [19:0] cfiType_20_pad;
  wire [13:0] cfiType_22_shl;
  wire [19:0] cfiType_22_pad;
  wire [13:0] cfiType_23_shl;
  wire [19:0] cfiType_23_pad;
  wire [13:0] cfiType_0_shl;
  wire [19:0] cfiType_0_pad;
  wire [9:0] tgtPages_11_shl;
  wire [19:0] tgtPages_11_pad;
  wire [13:0] cfiType_7_shl;
  wire [19:0] cfiType_7_pad;
  wire [13:0] cfiType_19_shl;
  wire [19:0] cfiType_19_pad;
  wire [13:0] cfiType_17_shl;
  wire [19:0] cfiType_17_pad;
  wire [13:0] cfiType_25_shl;
  wire [19:0] cfiType_25_pad;
  wire [13:0] cfiType_3_shl;
  wire [19:0] cfiType_3_pad;
  wire [13:0] cfiType_10_shl;
  wire [19:0] cfiType_10_pad;
  wire [9:0] tgtPages_14_shl;
  wire [19:0] tgtPages_14_pad;
  wire [13:0] cfiType_2_shl;
  wire [19:0] cfiType_2_pad;
  wire [13:0] cfiType_16_shl;
  wire [19:0] cfiType_16_pad;
  wire [9:0] tgtPages_0_shl;
  wire [19:0] tgtPages_0_pad;
  wire [9:0] tgtPages_21_shl;
  wire [19:0] tgtPages_21_pad;
  wire [9:0] tgtPages_5_shl;
  wire [19:0] tgtPages_5_pad;
  wire [9:0] tgtPages_4_shl;
  wire [19:0] tgtPages_4_pad;
  wire [13:0] cfiType_9_shl;
  wire [19:0] cfiType_9_pad;
  wire [9:0] tgtPages_25_shl;
  wire [19:0] tgtPages_25_pad;
  wire [13:0] cfiType_8_shl;
  wire [19:0] cfiType_8_pad;
  wire [9:0] tgtPages_24_shl;
  wire [19:0] tgtPages_24_pad;
  wire [13:0] cfiType_26_shl;
  wire [19:0] cfiType_26_pad;
  wire [9:0] tgtPages_13_shl;
  wire [19:0] tgtPages_13_pad;
  wire [13:0] cfiType_14_shl;
  wire [19:0] cfiType_14_pad;
  wire [13:0] cfiType_11_shl;
  wire [19:0] cfiType_11_pad;
  wire [9:0] tgtPages_16_shl;
  wire [19:0] tgtPages_16_pad;
  wire [13:0] cfiType_15_shl;
  wire [19:0] cfiType_15_pad;
  wire [13:0] cfiType_24_shl;
  wire [19:0] cfiType_24_pad;
  wire [9:0] tgtPages_18_shl;
  wire [19:0] tgtPages_18_pad;
  wire [13:0] cfiType_21_shl;
  wire [19:0] cfiType_21_pad;
  wire [9:0] tgtPages_12_shl;
  wire [19:0] tgtPages_12_pad;
  wire [9:0] tgtPages_10_shl;
  wire [19:0] tgtPages_10_pad;
  wire [9:0] tgtPages_15_shl;
  wire [19:0] tgtPages_15_pad;
  wire [9:0] tgtPages_22_shl;
  wire [19:0] tgtPages_22_pad;
  wire [9:0] tgtPages_19_shl;
  wire [19:0] tgtPages_19_pad;
  wire [13:0] cfiType_13_shl;
  wire [19:0] cfiType_13_pad;
  wire [13:0] cfiType_6_shl;
  wire [19:0] cfiType_6_pad;
  wire [9:0] tgtPages_6_shl;
  wire [19:0] tgtPages_6_pad;
  wire [13:0] cfiType_27_shl;
  wire [19:0] cfiType_27_pad;
  wire [9:0] tgtPages_23_shl;
  wire [19:0] tgtPages_23_pad;
  wire [13:0] cfiType_12_shl;
  wire [19:0] cfiType_12_pad;
  wire [9:0] tgtPages_8_shl;
  wire [19:0] tgtPages_8_pad;
  wire [9:0] tgtPages_1_shl;
  wire [19:0] tgtPages_1_pad;
  wire [9:0] tgtPages_9_shl;
  wire [19:0] tgtPages_9_pad;
  wire [13:0] cfiType_5_shl;
  wire [19:0] cfiType_5_pad;
  wire [9:0] tgtPages_7_shl;
  wire [19:0] tgtPages_7_pad;
  wire [9:0] tgtPages_27_shl;
  wire [19:0] tgtPages_27_pad;
  wire [19:0] BTB_xor31;
  wire [19:0] BTB_xor66;
  wire [19:0] BTB_xor32;
  wire [19:0] BTB_xor15;
  wire [19:0] BTB_xor68;
  wire [19:0] BTB_xor33;
  wire [19:0] BTB_xor70;
  wire [19:0] BTB_xor34;
  wire [19:0] BTB_xor16;
  wire [19:0] BTB_xor7;
  wire [19:0] BTB_xor72;
  wire [19:0] BTB_xor35;
  wire [19:0] BTB_xor74;
  wire [19:0] BTB_xor36;
  wire [19:0] BTB_xor17;
  wire [19:0] BTB_xor76;
  wire [19:0] BTB_xor37;
  wire [19:0] BTB_xor78;
  wire [19:0] BTB_xor38;
  wire [19:0] BTB_xor18;
  wire [19:0] BTB_xor8;
  wire [19:0] BTB_xor3;
  wire [19:0] BTB_xor39;
  wire [19:0] BTB_xor82;
  wire [19:0] BTB_xor40;
  wire [19:0] BTB_xor19;
  wire [19:0] BTB_xor84;
  wire [19:0] BTB_xor41;
  wire [19:0] BTB_xor86;
  wire [19:0] BTB_xor42;
  wire [19:0] BTB_xor20;
  wire [19:0] BTB_xor9;
  wire [19:0] BTB_xor88;
  wire [19:0] BTB_xor43;
  wire [19:0] BTB_xor90;
  wire [19:0] BTB_xor44;
  wire [19:0] BTB_xor21;
  wire [19:0] BTB_xor92;
  wire [19:0] BTB_xor45;
  wire [19:0] BTB_xor94;
  wire [19:0] BTB_xor46;
  wire [19:0] BTB_xor22;
  wire [19:0] BTB_xor10;
  wire [19:0] BTB_xor4;
  wire [19:0] BTB_xor1;
  wire [19:0] BTB_xor47;
  wire [19:0] BTB_xor98;
  wire [19:0] BTB_xor48;
  wire [19:0] BTB_xor23;
  wire [19:0] BTB_xor100;
  wire [19:0] BTB_xor49;
  wire [19:0] BTB_xor102;
  wire [19:0] BTB_xor50;
  wire [19:0] BTB_xor24;
  wire [19:0] BTB_xor11;
  wire [19:0] BTB_xor104;
  wire [19:0] BTB_xor51;
  wire [19:0] BTB_xor106;
  wire [19:0] BTB_xor52;
  wire [19:0] BTB_xor25;
  wire [19:0] BTB_xor108;
  wire [19:0] BTB_xor53;
  wire [19:0] BTB_xor110;
  wire [19:0] BTB_xor54;
  wire [19:0] BTB_xor26;
  wire [19:0] BTB_xor12;
  wire [19:0] BTB_xor5;
  wire [19:0] BTB_xor112;
  wire [19:0] BTB_xor55;
  wire [19:0] BTB_xor114;
  wire [19:0] BTB_xor56;
  wire [19:0] BTB_xor27;
  wire [19:0] BTB_xor116;
  wire [19:0] BTB_xor57;
  wire [19:0] BTB_xor118;
  wire [19:0] BTB_xor58;
  wire [19:0] BTB_xor28;
  wire [19:0] BTB_xor13;
  wire [19:0] BTB_xor120;
  wire [19:0] BTB_xor59;
  wire [19:0] BTB_xor122;
  wire [19:0] BTB_xor60;
  wire [19:0] BTB_xor29;
  wire [19:0] BTB_xor124;
  wire [19:0] BTB_xor61;
  wire [19:0] BTB_xor126;
  wire [19:0] BTB_xor62;
  wire [19:0] BTB_xor30;
  wire [19:0] BTB_xor14;
  wire [19:0] BTB_xor6;
  wire [19:0] BTB_xor2;
  wire [19:0] BTB_xor0;
  assign _T_1037__T_1106_addr = _T_1101 ^ _T_1104;
  assign _T_1037__T_1106_data = _T_1037[_T_1037__T_1106_addr]; // @[BTB.scala 113:26]
  assign _T_1037__T_1119_data = io_bht_update_bits_taken;
  assign _T_1037__T_1119_addr = _T_1114 ^ _T_1117;
  assign _T_1037__T_1119_mask = 1'h1;
  assign _T_1037__T_1119_en = io_bht_update_valid & io_bht_update_bits_branch;
  assign _T_1 = pages_0 == io_req_bits_addr[38:14]; // @[BTB.scala 202:29]
  assign _T_2 = pages_1 == io_req_bits_addr[38:14]; // @[BTB.scala 202:29]
  assign _T_3 = pages_2 == io_req_bits_addr[38:14]; // @[BTB.scala 202:29]
  assign _T_4 = pages_3 == io_req_bits_addr[38:14]; // @[BTB.scala 202:29]
  assign _T_5 = pages_4 == io_req_bits_addr[38:14]; // @[BTB.scala 202:29]
  assign _T_6 = pages_5 == io_req_bits_addr[38:14]; // @[BTB.scala 202:29]
  assign _T_11 = {_T_6,_T_5,_T_4,_T_3,_T_2,_T_1}; // @[Cat.scala 29:58]
  assign pageHit = pageValid & _T_11; // @[BTB.scala 202:15]
  assign _T_13 = idxs_0 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_14 = idxs_1 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_15 = idxs_2 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_16 = idxs_3 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_17 = idxs_4 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_18 = idxs_5 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_19 = idxs_6 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_20 = idxs_7 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_21 = idxs_8 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_22 = idxs_9 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_23 = idxs_10 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_24 = idxs_11 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_25 = idxs_12 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_26 = idxs_13 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_27 = idxs_14 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_28 = idxs_15 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_29 = idxs_16 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_30 = idxs_17 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_31 = idxs_18 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_32 = idxs_19 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_33 = idxs_20 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_34 = idxs_21 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_35 = idxs_22 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_36 = idxs_23 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_37 = idxs_24 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_38 = idxs_25 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_39 = idxs_26 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_40 = idxs_27 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_46 = {_T_19,_T_18,_T_17,_T_16,_T_15,_T_14,_T_13}; // @[Cat.scala 29:58]
  assign _T_53 = {_T_26,_T_25,_T_24,_T_23,_T_22,_T_21,_T_20,_T_46}; // @[Cat.scala 29:58]
  assign _T_59 = {_T_33,_T_32,_T_31,_T_30,_T_29,_T_28,_T_27}; // @[Cat.scala 29:58]
  assign _T_67 = {_T_40,_T_39,_T_38,_T_37,_T_36,_T_35,_T_34,_T_59,_T_53}; // @[Cat.scala 29:58]
  assign idxHit = _T_67 & isValid; // @[BTB.scala 206:32]
  assign _T_69 = pages_0 == r_btb_updatePipe_bits_pc[38:14]; // @[BTB.scala 202:29]
  assign _T_70 = pages_1 == r_btb_updatePipe_bits_pc[38:14]; // @[BTB.scala 202:29]
  assign _T_71 = pages_2 == r_btb_updatePipe_bits_pc[38:14]; // @[BTB.scala 202:29]
  assign _T_72 = pages_3 == r_btb_updatePipe_bits_pc[38:14]; // @[BTB.scala 202:29]
  assign _T_73 = pages_4 == r_btb_updatePipe_bits_pc[38:14]; // @[BTB.scala 202:29]
  assign _T_74 = pages_5 == r_btb_updatePipe_bits_pc[38:14]; // @[BTB.scala 202:29]
  assign _T_79 = {_T_74,_T_73,_T_72,_T_71,_T_70,_T_69}; // @[Cat.scala 29:58]
  assign updatePageHit = pageValid & _T_79; // @[BTB.scala 202:15]
  assign updateHit = r_btb_updatePipe_bits_prediction_entry < 5'h1c; // @[BTB.scala 220:48]
  assign useUpdatePageHit = |updatePageHit; // @[BTB.scala 222:40]
  assign usePageHit = |pageHit; // @[BTB.scala 223:28]
  assign doIdxPageRepl = ~useUpdatePageHit; // @[BTB.scala 224:23]
  assign _T_82 = {pageHit[4:0],pageHit[5]}; // @[Cat.scala 29:58]
  assign _T_83 = 8'h1 << nextPageRepl; // @[OneHot.scala 58:35]
  assign _T_84 = usePageHit ? 8'h0 : _T_83; // @[BTB.scala 226:70]
  assign _GEN_432 = {{2'd0}, _T_82}; // @[BTB.scala 226:65]
  assign idxPageRepl = _GEN_432 | _T_84; // @[BTB.scala 226:65]
  assign idxPageUpdateOH = useUpdatePageHit ? {{2'd0}, updatePageHit} : idxPageRepl; // @[BTB.scala 227:28]
  assign _T_87 = |idxPageUpdateOH[7:4]; // @[OneHot.scala 32:14]
  assign _T_88 = idxPageUpdateOH[7:4] | idxPageUpdateOH[3:0]; // @[OneHot.scala 32:28]
  assign _T_91 = |_T_88[3:2]; // @[OneHot.scala 32:14]
  assign _T_92 = _T_88[3:2] | _T_88[1:0]; // @[OneHot.scala 32:28]
  assign idxPageUpdate = {_T_87,_T_91,_T_92[1]}; // @[Cat.scala 29:58]
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 8'h0; // @[BTB.scala 229:26]
  assign samePage = r_btb_updatePipe_bits_pc[38:14] == io_req_bits_addr[38:14]; // @[BTB.scala 231:45]
  assign doTgtPageRepl = ~samePage & ~usePageHit; // @[BTB.scala 232:33]
  assign _T_101 = {idxPageUpdateOH[4:0],idxPageUpdateOH[5]}; // @[Cat.scala 29:58]
  assign tgtPageRepl = samePage ? idxPageUpdateOH : {{2'd0}, _T_101}; // @[BTB.scala 233:24]
  assign _T_102 = usePageHit ? 8'h0 : tgtPageRepl; // @[BTB.scala 234:45]
  assign _GEN_433 = {{2'd0}, pageHit}; // @[BTB.scala 234:40]
  assign _T_103 = _GEN_433 | _T_102; // @[BTB.scala 234:40]
  assign _T_106 = |_T_103[7:4]; // @[OneHot.scala 32:14]
  assign _T_107 = _T_103[7:4] | _T_103[3:0]; // @[OneHot.scala 32:28]
  assign _T_110 = |_T_107[3:2]; // @[OneHot.scala 32:14]
  assign _T_111 = _T_107[3:2] | _T_107[1:0]; // @[OneHot.scala 32:28]
  assign tgtPageUpdate = {_T_106,_T_110,_T_111[1]}; // @[Cat.scala 29:58]
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 8'h0; // @[BTB.scala 235:26]
  assign _T_114 = doIdxPageRepl | doTgtPageRepl; // @[BTB.scala 237:46]
  assign _T_115 = r_btb_updatePipe_valid & _T_114; // @[BTB.scala 237:28]
  assign _T_116 = doIdxPageRepl & doTgtPageRepl; // @[BTB.scala 238:30]
  assign _T_117 = _T_116 ? 2'h2 : 2'h1; // @[BTB.scala 239:40]
  assign _GEN_434 = {{1'd0}, _T_117}; // @[BTB.scala 239:29]
  assign _T_119 = nextPageRepl + _GEN_434; // @[BTB.scala 239:29]
  assign _T_120 = _T_119 >= 3'h6; // @[BTB.scala 240:30]
  assign _T_135 = _T_123[24] ? _T_123[23] : _T_123[22]; // @[Replacement.scala 240:16]
  assign _T_136 = {_T_123[24],_T_135}; // @[Cat.scala 29:58]
  assign _T_145 = _T_123[20] ? _T_123[19] : _T_123[18]; // @[Replacement.scala 240:16]
  assign _T_146 = {_T_123[20],_T_145}; // @[Cat.scala 29:58]
  assign _T_152 = _T_123[17] ? _T_123[16] : _T_123[15]; // @[Replacement.scala 240:16]
  assign _T_153 = {_T_123[17],_T_152}; // @[Cat.scala 29:58]
  assign _T_154 = _T_123[21] ? _T_146 : _T_153; // @[Replacement.scala 240:16]
  assign _T_155 = {_T_123[21],_T_154}; // @[Cat.scala 29:58]
  assign _T_156 = _T_123[25] ? {{1'd0}, _T_136} : _T_155; // @[Replacement.scala 240:16]
  assign _T_157 = {_T_123[25],_T_156}; // @[Cat.scala 29:58]
  assign _T_169 = _T_123[12] ? _T_123[11] : _T_123[10]; // @[Replacement.scala 240:16]
  assign _T_170 = {_T_123[12],_T_169}; // @[Cat.scala 29:58]
  assign _T_176 = _T_123[9] ? _T_123[8] : _T_123[7]; // @[Replacement.scala 240:16]
  assign _T_177 = {_T_123[9],_T_176}; // @[Cat.scala 29:58]
  assign _T_178 = _T_123[13] ? _T_170 : _T_177; // @[Replacement.scala 240:16]
  assign _T_179 = {_T_123[13],_T_178}; // @[Cat.scala 29:58]
  assign _T_188 = _T_123[5] ? _T_123[4] : _T_123[3]; // @[Replacement.scala 240:16]
  assign _T_189 = {_T_123[5],_T_188}; // @[Cat.scala 29:58]
  assign _T_195 = _T_123[2] ? _T_123[1] : _T_123[0]; // @[Replacement.scala 240:16]
  assign _T_196 = {_T_123[2],_T_195}; // @[Cat.scala 29:58]
  assign _T_197 = _T_123[6] ? _T_189 : _T_196; // @[Replacement.scala 240:16]
  assign _T_198 = {_T_123[6],_T_197}; // @[Cat.scala 29:58]
  assign _T_199 = _T_123[14] ? _T_179 : _T_198; // @[Replacement.scala 240:16]
  assign _T_200 = {_T_123[14],_T_199}; // @[Cat.scala 29:58]
  assign _T_201 = _T_123[26] ? _T_157 : _T_200; // @[Replacement.scala 240:16]
  assign _T_202 = {_T_123[26],_T_201}; // @[Cat.scala 29:58]
  assign waddr = updateHit ? r_btb_updatePipe_bits_prediction_entry : _T_202; // @[BTB.scala 244:18]
  assign _T_203 = r_respPipe_valid & r_respPipe_bits_taken; // @[BTB.scala 246:22]
  assign _T_204 = _T_203 | r_btb_updatePipe_valid; // @[BTB.scala 246:43]
  assign _T_205 = r_btb_updatePipe_valid ? waddr : r_respPipe_bits_entry; // @[BTB.scala 247:20]
  assign _T_224 = _T_205[1] ? ~_T_205[0] : _T_123[23]; // @[Replacement.scala 193:16]
  assign _T_228 = _T_205[1] ? _T_123[22] : ~_T_205[0]; // @[Replacement.scala 196:16]
  assign _T_230 = {~_T_205[1],_T_224,_T_228}; // @[Cat.scala 29:58]
  assign _T_231 = _T_205[3] ? _T_230 : _T_123[24:22]; // @[Replacement.scala 193:16]
  assign _T_245 = _T_205[1] ? ~_T_205[0] : _T_123[19]; // @[Replacement.scala 193:16]
  assign _T_249 = _T_205[1] ? _T_123[18] : ~_T_205[0]; // @[Replacement.scala 196:16]
  assign _T_251 = {~_T_205[1],_T_245,_T_249}; // @[Cat.scala 29:58]
  assign _T_252 = _T_205[2] ? _T_251 : _T_123[20:18]; // @[Replacement.scala 193:16]
  assign _T_261 = _T_205[1] ? ~_T_205[0] : _T_123[16]; // @[Replacement.scala 193:16]
  assign _T_265 = _T_205[1] ? _T_123[15] : ~_T_205[0]; // @[Replacement.scala 196:16]
  assign _T_267 = {~_T_205[1],_T_261,_T_265}; // @[Cat.scala 29:58]
  assign _T_268 = _T_205[2] ? _T_123[17:15] : _T_267; // @[Replacement.scala 196:16]
  assign _T_270 = {~_T_205[2],_T_252,_T_268}; // @[Cat.scala 29:58]
  assign _T_271 = _T_205[3] ? _T_123[21:15] : _T_270; // @[Replacement.scala 196:16]
  assign _T_273 = {~_T_205[3],_T_231,_T_271}; // @[Cat.scala 29:58]
  assign _T_274 = _T_205[4] ? _T_273 : _T_123[25:15]; // @[Replacement.scala 193:16]
  assign _T_293 = _T_205[1] ? ~_T_205[0] : _T_123[11]; // @[Replacement.scala 193:16]
  assign _T_297 = _T_205[1] ? _T_123[10] : ~_T_205[0]; // @[Replacement.scala 196:16]
  assign _T_299 = {~_T_205[1],_T_293,_T_297}; // @[Cat.scala 29:58]
  assign _T_300 = _T_205[2] ? _T_299 : _T_123[12:10]; // @[Replacement.scala 193:16]
  assign _T_309 = _T_205[1] ? ~_T_205[0] : _T_123[8]; // @[Replacement.scala 193:16]
  assign _T_313 = _T_205[1] ? _T_123[7] : ~_T_205[0]; // @[Replacement.scala 196:16]
  assign _T_315 = {~_T_205[1],_T_309,_T_313}; // @[Cat.scala 29:58]
  assign _T_316 = _T_205[2] ? _T_123[9:7] : _T_315; // @[Replacement.scala 196:16]
  assign _T_318 = {~_T_205[2],_T_300,_T_316}; // @[Cat.scala 29:58]
  assign _T_319 = _T_205[3] ? _T_318 : _T_123[13:7]; // @[Replacement.scala 193:16]
  assign _T_333 = _T_205[1] ? ~_T_205[0] : _T_123[4]; // @[Replacement.scala 193:16]
  assign _T_337 = _T_205[1] ? _T_123[3] : ~_T_205[0]; // @[Replacement.scala 196:16]
  assign _T_339 = {~_T_205[1],_T_333,_T_337}; // @[Cat.scala 29:58]
  assign _T_340 = _T_205[2] ? _T_339 : _T_123[5:3]; // @[Replacement.scala 193:16]
  assign _T_349 = _T_205[1] ? ~_T_205[0] : _T_123[1]; // @[Replacement.scala 193:16]
  assign _T_353 = _T_205[1] ? _T_123[0] : ~_T_205[0]; // @[Replacement.scala 196:16]
  assign _T_355 = {~_T_205[1],_T_349,_T_353}; // @[Cat.scala 29:58]
  assign _T_356 = _T_205[2] ? _T_123[2:0] : _T_355; // @[Replacement.scala 196:16]
  assign _T_358 = {~_T_205[2],_T_340,_T_356}; // @[Cat.scala 29:58]
  assign _T_359 = _T_205[3] ? _T_123[6:0] : _T_358; // @[Replacement.scala 196:16]
  assign _T_361 = {~_T_205[3],_T_319,_T_359}; // @[Cat.scala 29:58]
  assign _T_362 = _T_205[4] ? _T_123[14:0] : _T_361; // @[Replacement.scala 196:16]
  assign _T_364 = {~_T_205[4],_T_274,_T_362}; // @[Cat.scala 29:58]
  assign _T_365 = 32'h1 << waddr; // @[OneHot.scala 58:35]
  assign _T_368 = idxPageUpdate + 3'h1; // @[BTB.scala 254:38]
  assign _GEN_435 = {{4'd0}, isValid}; // @[BTB.scala 257:55]
  assign _T_369 = _GEN_435 | _T_365; // @[BTB.scala 257:55]
  assign _T_371 = _GEN_435 & ~_T_365; // @[BTB.scala 257:71]
  assign _T_372 = r_btb_updatePipe_bits_isValid ? _T_369 : _T_371; // @[BTB.scala 257:19]
  assign _T_376 = idxPageUpdate[0] ? tgtPageReplEn : idxPageReplEn; // @[BTB.scala 268:24]
  assign _T_383 = idxPageUpdate[0] ? idxPageReplEn : tgtPageReplEn; // @[BTB.scala 270:24]
  assign _GEN_437 = {{2'd0}, pageValid}; // @[BTB.scala 272:28]
  assign _T_390 = _GEN_437 | tgtPageReplEn; // @[BTB.scala 272:28]
  assign _T_391 = _T_390 | idxPageReplEn; // @[BTB.scala 272:44]
  assign _GEN_338 = r_btb_updatePipe_valid ? _T_372 : {{4'd0}, isValid}; // @[BTB.scala 250:29]
  assign _GEN_373 = r_btb_updatePipe_valid ? _T_391 : {{2'd0}, pageValid}; // @[BTB.scala 250:29]
  assign _T_392 = {pageHit, 1'h0}; // @[BTB.scala 275:29]
  assign _T_421 = idxHit[0] ? idxPages_0 : 3'h0; // @[Mux.scala 27:72]
  assign _T_422 = idxHit[1] ? idxPages_1 : 3'h0; // @[Mux.scala 27:72]
  assign _T_423 = idxHit[2] ? idxPages_2 : 3'h0; // @[Mux.scala 27:72]
  assign _T_424 = idxHit[3] ? idxPages_3 : 3'h0; // @[Mux.scala 27:72]
  assign _T_425 = idxHit[4] ? idxPages_4 : 3'h0; // @[Mux.scala 27:72]
  assign _T_426 = idxHit[5] ? idxPages_5 : 3'h0; // @[Mux.scala 27:72]
  assign _T_427 = idxHit[6] ? idxPages_6 : 3'h0; // @[Mux.scala 27:72]
  assign _T_428 = idxHit[7] ? idxPages_7 : 3'h0; // @[Mux.scala 27:72]
  assign _T_429 = idxHit[8] ? idxPages_8 : 3'h0; // @[Mux.scala 27:72]
  assign _T_430 = idxHit[9] ? idxPages_9 : 3'h0; // @[Mux.scala 27:72]
  assign _T_431 = idxHit[10] ? idxPages_10 : 3'h0; // @[Mux.scala 27:72]
  assign _T_432 = idxHit[11] ? idxPages_11 : 3'h0; // @[Mux.scala 27:72]
  assign _T_433 = idxHit[12] ? idxPages_12 : 3'h0; // @[Mux.scala 27:72]
  assign _T_434 = idxHit[13] ? idxPages_13 : 3'h0; // @[Mux.scala 27:72]
  assign _T_435 = idxHit[14] ? idxPages_14 : 3'h0; // @[Mux.scala 27:72]
  assign _T_436 = idxHit[15] ? idxPages_15 : 3'h0; // @[Mux.scala 27:72]
  assign _T_437 = idxHit[16] ? idxPages_16 : 3'h0; // @[Mux.scala 27:72]
  assign _T_438 = idxHit[17] ? idxPages_17 : 3'h0; // @[Mux.scala 27:72]
  assign _T_439 = idxHit[18] ? idxPages_18 : 3'h0; // @[Mux.scala 27:72]
  assign _T_440 = idxHit[19] ? idxPages_19 : 3'h0; // @[Mux.scala 27:72]
  assign _T_441 = idxHit[20] ? idxPages_20 : 3'h0; // @[Mux.scala 27:72]
  assign _T_442 = idxHit[21] ? idxPages_21 : 3'h0; // @[Mux.scala 27:72]
  assign _T_443 = idxHit[22] ? idxPages_22 : 3'h0; // @[Mux.scala 27:72]
  assign _T_444 = idxHit[23] ? idxPages_23 : 3'h0; // @[Mux.scala 27:72]
  assign _T_445 = idxHit[24] ? idxPages_24 : 3'h0; // @[Mux.scala 27:72]
  assign _T_446 = idxHit[25] ? idxPages_25 : 3'h0; // @[Mux.scala 27:72]
  assign _T_447 = idxHit[26] ? idxPages_26 : 3'h0; // @[Mux.scala 27:72]
  assign _T_448 = idxHit[27] ? idxPages_27 : 3'h0; // @[Mux.scala 27:72]
  assign _T_449 = _T_421 | _T_422; // @[Mux.scala 27:72]
  assign _T_450 = _T_449 | _T_423; // @[Mux.scala 27:72]
  assign _T_451 = _T_450 | _T_424; // @[Mux.scala 27:72]
  assign _T_452 = _T_451 | _T_425; // @[Mux.scala 27:72]
  assign _T_453 = _T_452 | _T_426; // @[Mux.scala 27:72]
  assign _T_454 = _T_453 | _T_427; // @[Mux.scala 27:72]
  assign _T_455 = _T_454 | _T_428; // @[Mux.scala 27:72]
  assign _T_456 = _T_455 | _T_429; // @[Mux.scala 27:72]
  assign _T_457 = _T_456 | _T_430; // @[Mux.scala 27:72]
  assign _T_458 = _T_457 | _T_431; // @[Mux.scala 27:72]
  assign _T_459 = _T_458 | _T_432; // @[Mux.scala 27:72]
  assign _T_460 = _T_459 | _T_433; // @[Mux.scala 27:72]
  assign _T_461 = _T_460 | _T_434; // @[Mux.scala 27:72]
  assign _T_462 = _T_461 | _T_435; // @[Mux.scala 27:72]
  assign _T_463 = _T_462 | _T_436; // @[Mux.scala 27:72]
  assign _T_464 = _T_463 | _T_437; // @[Mux.scala 27:72]
  assign _T_465 = _T_464 | _T_438; // @[Mux.scala 27:72]
  assign _T_466 = _T_465 | _T_439; // @[Mux.scala 27:72]
  assign _T_467 = _T_466 | _T_440; // @[Mux.scala 27:72]
  assign _T_468 = _T_467 | _T_441; // @[Mux.scala 27:72]
  assign _T_469 = _T_468 | _T_442; // @[Mux.scala 27:72]
  assign _T_470 = _T_469 | _T_443; // @[Mux.scala 27:72]
  assign _T_471 = _T_470 | _T_444; // @[Mux.scala 27:72]
  assign _T_472 = _T_471 | _T_445; // @[Mux.scala 27:72]
  assign _T_473 = _T_472 | _T_446; // @[Mux.scala 27:72]
  assign _T_474 = _T_473 | _T_447; // @[Mux.scala 27:72]
  assign _T_475 = _T_474 | _T_448; // @[Mux.scala 27:72]
  assign _T_477 = _T_392 >> _T_475; // @[BTB.scala 275:34]
  assign _T_507 = idxHit[0] ? tgtPages_0 : 3'h0; // @[Mux.scala 27:72]
  assign _T_508 = idxHit[1] ? tgtPages_1 : 3'h0; // @[Mux.scala 27:72]
  assign _T_509 = idxHit[2] ? tgtPages_2 : 3'h0; // @[Mux.scala 27:72]
  assign _T_510 = idxHit[3] ? tgtPages_3 : 3'h0; // @[Mux.scala 27:72]
  assign _T_511 = idxHit[4] ? tgtPages_4 : 3'h0; // @[Mux.scala 27:72]
  assign _T_512 = idxHit[5] ? tgtPages_5 : 3'h0; // @[Mux.scala 27:72]
  assign _T_513 = idxHit[6] ? tgtPages_6 : 3'h0; // @[Mux.scala 27:72]
  assign _T_514 = idxHit[7] ? tgtPages_7 : 3'h0; // @[Mux.scala 27:72]
  assign _T_515 = idxHit[8] ? tgtPages_8 : 3'h0; // @[Mux.scala 27:72]
  assign _T_516 = idxHit[9] ? tgtPages_9 : 3'h0; // @[Mux.scala 27:72]
  assign _T_517 = idxHit[10] ? tgtPages_10 : 3'h0; // @[Mux.scala 27:72]
  assign _T_518 = idxHit[11] ? tgtPages_11 : 3'h0; // @[Mux.scala 27:72]
  assign _T_519 = idxHit[12] ? tgtPages_12 : 3'h0; // @[Mux.scala 27:72]
  assign _T_520 = idxHit[13] ? tgtPages_13 : 3'h0; // @[Mux.scala 27:72]
  assign _T_521 = idxHit[14] ? tgtPages_14 : 3'h0; // @[Mux.scala 27:72]
  assign _T_522 = idxHit[15] ? tgtPages_15 : 3'h0; // @[Mux.scala 27:72]
  assign _T_523 = idxHit[16] ? tgtPages_16 : 3'h0; // @[Mux.scala 27:72]
  assign _T_524 = idxHit[17] ? tgtPages_17 : 3'h0; // @[Mux.scala 27:72]
  assign _T_525 = idxHit[18] ? tgtPages_18 : 3'h0; // @[Mux.scala 27:72]
  assign _T_526 = idxHit[19] ? tgtPages_19 : 3'h0; // @[Mux.scala 27:72]
  assign _T_527 = idxHit[20] ? tgtPages_20 : 3'h0; // @[Mux.scala 27:72]
  assign _T_528 = idxHit[21] ? tgtPages_21 : 3'h0; // @[Mux.scala 27:72]
  assign _T_529 = idxHit[22] ? tgtPages_22 : 3'h0; // @[Mux.scala 27:72]
  assign _T_530 = idxHit[23] ? tgtPages_23 : 3'h0; // @[Mux.scala 27:72]
  assign _T_531 = idxHit[24] ? tgtPages_24 : 3'h0; // @[Mux.scala 27:72]
  assign _T_532 = idxHit[25] ? tgtPages_25 : 3'h0; // @[Mux.scala 27:72]
  assign _T_533 = idxHit[26] ? tgtPages_26 : 3'h0; // @[Mux.scala 27:72]
  assign _T_534 = idxHit[27] ? tgtPages_27 : 3'h0; // @[Mux.scala 27:72]
  assign _T_535 = _T_507 | _T_508; // @[Mux.scala 27:72]
  assign _T_536 = _T_535 | _T_509; // @[Mux.scala 27:72]
  assign _T_537 = _T_536 | _T_510; // @[Mux.scala 27:72]
  assign _T_538 = _T_537 | _T_511; // @[Mux.scala 27:72]
  assign _T_539 = _T_538 | _T_512; // @[Mux.scala 27:72]
  assign _T_540 = _T_539 | _T_513; // @[Mux.scala 27:72]
  assign _T_541 = _T_540 | _T_514; // @[Mux.scala 27:72]
  assign _T_542 = _T_541 | _T_515; // @[Mux.scala 27:72]
  assign _T_543 = _T_542 | _T_516; // @[Mux.scala 27:72]
  assign _T_544 = _T_543 | _T_517; // @[Mux.scala 27:72]
  assign _T_545 = _T_544 | _T_518; // @[Mux.scala 27:72]
  assign _T_546 = _T_545 | _T_519; // @[Mux.scala 27:72]
  assign _T_547 = _T_546 | _T_520; // @[Mux.scala 27:72]
  assign _T_548 = _T_547 | _T_521; // @[Mux.scala 27:72]
  assign _T_549 = _T_548 | _T_522; // @[Mux.scala 27:72]
  assign _T_550 = _T_549 | _T_523; // @[Mux.scala 27:72]
  assign _T_551 = _T_550 | _T_524; // @[Mux.scala 27:72]
  assign _T_552 = _T_551 | _T_525; // @[Mux.scala 27:72]
  assign _T_553 = _T_552 | _T_526; // @[Mux.scala 27:72]
  assign _T_554 = _T_553 | _T_527; // @[Mux.scala 27:72]
  assign _T_555 = _T_554 | _T_528; // @[Mux.scala 27:72]
  assign _T_556 = _T_555 | _T_529; // @[Mux.scala 27:72]
  assign _T_557 = _T_556 | _T_530; // @[Mux.scala 27:72]
  assign _T_558 = _T_557 | _T_531; // @[Mux.scala 27:72]
  assign _T_559 = _T_558 | _T_532; // @[Mux.scala 27:72]
  assign _T_560 = _T_559 | _T_533; // @[Mux.scala 27:72]
  assign _T_561 = _T_560 | _T_534; // @[Mux.scala 27:72]
  assign _T_591 = idxHit[0] ? tgts_0 : 13'h0; // @[Mux.scala 27:72]
  assign _T_592 = idxHit[1] ? tgts_1 : 13'h0; // @[Mux.scala 27:72]
  assign _T_593 = idxHit[2] ? tgts_2 : 13'h0; // @[Mux.scala 27:72]
  assign _T_594 = idxHit[3] ? tgts_3 : 13'h0; // @[Mux.scala 27:72]
  assign _T_595 = idxHit[4] ? tgts_4 : 13'h0; // @[Mux.scala 27:72]
  assign _T_596 = idxHit[5] ? tgts_5 : 13'h0; // @[Mux.scala 27:72]
  assign _T_597 = idxHit[6] ? tgts_6 : 13'h0; // @[Mux.scala 27:72]
  assign _T_598 = idxHit[7] ? tgts_7 : 13'h0; // @[Mux.scala 27:72]
  assign _T_599 = idxHit[8] ? tgts_8 : 13'h0; // @[Mux.scala 27:72]
  assign _T_600 = idxHit[9] ? tgts_9 : 13'h0; // @[Mux.scala 27:72]
  assign _T_601 = idxHit[10] ? tgts_10 : 13'h0; // @[Mux.scala 27:72]
  assign _T_602 = idxHit[11] ? tgts_11 : 13'h0; // @[Mux.scala 27:72]
  assign _T_603 = idxHit[12] ? tgts_12 : 13'h0; // @[Mux.scala 27:72]
  assign _T_604 = idxHit[13] ? tgts_13 : 13'h0; // @[Mux.scala 27:72]
  assign _T_605 = idxHit[14] ? tgts_14 : 13'h0; // @[Mux.scala 27:72]
  assign _T_606 = idxHit[15] ? tgts_15 : 13'h0; // @[Mux.scala 27:72]
  assign _T_607 = idxHit[16] ? tgts_16 : 13'h0; // @[Mux.scala 27:72]
  assign _T_608 = idxHit[17] ? tgts_17 : 13'h0; // @[Mux.scala 27:72]
  assign _T_609 = idxHit[18] ? tgts_18 : 13'h0; // @[Mux.scala 27:72]
  assign _T_610 = idxHit[19] ? tgts_19 : 13'h0; // @[Mux.scala 27:72]
  assign _T_611 = idxHit[20] ? tgts_20 : 13'h0; // @[Mux.scala 27:72]
  assign _T_612 = idxHit[21] ? tgts_21 : 13'h0; // @[Mux.scala 27:72]
  assign _T_613 = idxHit[22] ? tgts_22 : 13'h0; // @[Mux.scala 27:72]
  assign _T_614 = idxHit[23] ? tgts_23 : 13'h0; // @[Mux.scala 27:72]
  assign _T_615 = idxHit[24] ? tgts_24 : 13'h0; // @[Mux.scala 27:72]
  assign _T_616 = idxHit[25] ? tgts_25 : 13'h0; // @[Mux.scala 27:72]
  assign _T_617 = idxHit[26] ? tgts_26 : 13'h0; // @[Mux.scala 27:72]
  assign _T_618 = idxHit[27] ? tgts_27 : 13'h0; // @[Mux.scala 27:72]
  assign _T_619 = _T_591 | _T_592; // @[Mux.scala 27:72]
  assign _T_620 = _T_619 | _T_593; // @[Mux.scala 27:72]
  assign _T_621 = _T_620 | _T_594; // @[Mux.scala 27:72]
  assign _T_622 = _T_621 | _T_595; // @[Mux.scala 27:72]
  assign _T_623 = _T_622 | _T_596; // @[Mux.scala 27:72]
  assign _T_624 = _T_623 | _T_597; // @[Mux.scala 27:72]
  assign _T_625 = _T_624 | _T_598; // @[Mux.scala 27:72]
  assign _T_626 = _T_625 | _T_599; // @[Mux.scala 27:72]
  assign _T_627 = _T_626 | _T_600; // @[Mux.scala 27:72]
  assign _T_628 = _T_627 | _T_601; // @[Mux.scala 27:72]
  assign _T_629 = _T_628 | _T_602; // @[Mux.scala 27:72]
  assign _T_630 = _T_629 | _T_603; // @[Mux.scala 27:72]
  assign _T_631 = _T_630 | _T_604; // @[Mux.scala 27:72]
  assign _T_632 = _T_631 | _T_605; // @[Mux.scala 27:72]
  assign _T_633 = _T_632 | _T_606; // @[Mux.scala 27:72]
  assign _T_634 = _T_633 | _T_607; // @[Mux.scala 27:72]
  assign _T_635 = _T_634 | _T_608; // @[Mux.scala 27:72]
  assign _T_636 = _T_635 | _T_609; // @[Mux.scala 27:72]
  assign _T_637 = _T_636 | _T_610; // @[Mux.scala 27:72]
  assign _T_638 = _T_637 | _T_611; // @[Mux.scala 27:72]
  assign _T_639 = _T_638 | _T_612; // @[Mux.scala 27:72]
  assign _T_640 = _T_639 | _T_613; // @[Mux.scala 27:72]
  assign _T_641 = _T_640 | _T_614; // @[Mux.scala 27:72]
  assign _T_642 = _T_641 | _T_615; // @[Mux.scala 27:72]
  assign _T_643 = _T_642 | _T_616; // @[Mux.scala 27:72]
  assign _T_644 = _T_643 | _T_617; // @[Mux.scala 27:72]
  assign _T_645 = _T_644 | _T_618; // @[Mux.scala 27:72]
  assign _T_647 = {_T_645, 1'h0}; // @[BTB.scala 277:82]
  assign _GEN_375 = 3'h1 == _T_561 ? pages_1 : pages_0; // @[Cat.scala 29:58]
  assign _GEN_376 = 3'h2 == _T_561 ? pages_2 : _GEN_375; // @[Cat.scala 29:58]
  assign _GEN_377 = 3'h3 == _T_561 ? pages_3 : _GEN_376; // @[Cat.scala 29:58]
  assign _GEN_378 = 3'h4 == _T_561 ? pages_4 : _GEN_377; // @[Cat.scala 29:58]
  assign _GEN_379 = 3'h5 == _T_561 ? pages_5 : _GEN_378; // @[Cat.scala 29:58]
  assign _T_648 = {_GEN_379,_T_647}; // @[Cat.scala 29:58]
  assign _T_651 = |idxHit[27:16]; // @[OneHot.scala 32:14]
  assign _GEN_438 = {{4'd0}, idxHit[27:16]}; // @[OneHot.scala 32:28]
  assign _T_652 = _GEN_438 | idxHit[15:0]; // @[OneHot.scala 32:28]
  assign _T_655 = |_T_652[15:8]; // @[OneHot.scala 32:14]
  assign _T_656 = _T_652[15:8] | _T_652[7:0]; // @[OneHot.scala 32:28]
  assign _T_659 = |_T_656[7:4]; // @[OneHot.scala 32:14]
  assign _T_660 = _T_656[7:4] | _T_656[3:0]; // @[OneHot.scala 32:28]
  assign _T_663 = |_T_660[3:2]; // @[OneHot.scala 32:14]
  assign _T_664 = _T_660[3:2] | _T_660[1:0]; // @[OneHot.scala 32:28]
  assign _T_668 = {_T_655,_T_659,_T_663,_T_664[1]}; // @[Cat.scala 29:58]
  assign _T_698 = idxHit[0] & brIdx_0; // @[Mux.scala 27:72]
  assign _T_699 = idxHit[1] & brIdx_1; // @[Mux.scala 27:72]
  assign _T_700 = idxHit[2] & brIdx_2; // @[Mux.scala 27:72]
  assign _T_701 = idxHit[3] & brIdx_3; // @[Mux.scala 27:72]
  assign _T_702 = idxHit[4] & brIdx_4; // @[Mux.scala 27:72]
  assign _T_703 = idxHit[5] & brIdx_5; // @[Mux.scala 27:72]
  assign _T_704 = idxHit[6] & brIdx_6; // @[Mux.scala 27:72]
  assign _T_705 = idxHit[7] & brIdx_7; // @[Mux.scala 27:72]
  assign _T_706 = idxHit[8] & brIdx_8; // @[Mux.scala 27:72]
  assign _T_707 = idxHit[9] & brIdx_9; // @[Mux.scala 27:72]
  assign _T_708 = idxHit[10] & brIdx_10; // @[Mux.scala 27:72]
  assign _T_709 = idxHit[11] & brIdx_11; // @[Mux.scala 27:72]
  assign _T_710 = idxHit[12] & brIdx_12; // @[Mux.scala 27:72]
  assign _T_711 = idxHit[13] & brIdx_13; // @[Mux.scala 27:72]
  assign _T_712 = idxHit[14] & brIdx_14; // @[Mux.scala 27:72]
  assign _T_713 = idxHit[15] & brIdx_15; // @[Mux.scala 27:72]
  assign _T_714 = idxHit[16] & brIdx_16; // @[Mux.scala 27:72]
  assign _T_715 = idxHit[17] & brIdx_17; // @[Mux.scala 27:72]
  assign _T_716 = idxHit[18] & brIdx_18; // @[Mux.scala 27:72]
  assign _T_717 = idxHit[19] & brIdx_19; // @[Mux.scala 27:72]
  assign _T_718 = idxHit[20] & brIdx_20; // @[Mux.scala 27:72]
  assign _T_719 = idxHit[21] & brIdx_21; // @[Mux.scala 27:72]
  assign _T_720 = idxHit[22] & brIdx_22; // @[Mux.scala 27:72]
  assign _T_721 = idxHit[23] & brIdx_23; // @[Mux.scala 27:72]
  assign _T_722 = idxHit[24] & brIdx_24; // @[Mux.scala 27:72]
  assign _T_723 = idxHit[25] & brIdx_25; // @[Mux.scala 27:72]
  assign _T_724 = idxHit[26] & brIdx_26; // @[Mux.scala 27:72]
  assign _T_725 = idxHit[27] & brIdx_27; // @[Mux.scala 27:72]
  assign _T_726 = _T_698 | _T_699; // @[Mux.scala 27:72]
  assign _T_727 = _T_726 | _T_700; // @[Mux.scala 27:72]
  assign _T_728 = _T_727 | _T_701; // @[Mux.scala 27:72]
  assign _T_729 = _T_728 | _T_702; // @[Mux.scala 27:72]
  assign _T_730 = _T_729 | _T_703; // @[Mux.scala 27:72]
  assign _T_731 = _T_730 | _T_704; // @[Mux.scala 27:72]
  assign _T_732 = _T_731 | _T_705; // @[Mux.scala 27:72]
  assign _T_733 = _T_732 | _T_706; // @[Mux.scala 27:72]
  assign _T_734 = _T_733 | _T_707; // @[Mux.scala 27:72]
  assign _T_735 = _T_734 | _T_708; // @[Mux.scala 27:72]
  assign _T_736 = _T_735 | _T_709; // @[Mux.scala 27:72]
  assign _T_737 = _T_736 | _T_710; // @[Mux.scala 27:72]
  assign _T_738 = _T_737 | _T_711; // @[Mux.scala 27:72]
  assign _T_739 = _T_738 | _T_712; // @[Mux.scala 27:72]
  assign _T_740 = _T_739 | _T_713; // @[Mux.scala 27:72]
  assign _T_741 = _T_740 | _T_714; // @[Mux.scala 27:72]
  assign _T_742 = _T_741 | _T_715; // @[Mux.scala 27:72]
  assign _T_743 = _T_742 | _T_716; // @[Mux.scala 27:72]
  assign _T_744 = _T_743 | _T_717; // @[Mux.scala 27:72]
  assign _T_745 = _T_744 | _T_718; // @[Mux.scala 27:72]
  assign _T_746 = _T_745 | _T_719; // @[Mux.scala 27:72]
  assign _T_747 = _T_746 | _T_720; // @[Mux.scala 27:72]
  assign _T_748 = _T_747 | _T_721; // @[Mux.scala 27:72]
  assign _T_749 = _T_748 | _T_722; // @[Mux.scala 27:72]
  assign _T_750 = _T_749 | _T_723; // @[Mux.scala 27:72]
  assign _T_751 = _T_750 | _T_724; // @[Mux.scala 27:72]
  assign _T_855 = idxHit[1] | idxHit[2]; // @[Misc.scala 182:16]
  assign _T_857 = idxHit[1] & idxHit[2]; // @[Misc.scala 182:61]
  assign _T_859 = idxHit[0] | _T_855; // @[Misc.scala 182:16]
  assign _T_861 = idxHit[0] & _T_855; // @[Misc.scala 182:61]
  assign _T_862 = _T_857 | _T_861; // @[Misc.scala 182:49]
  assign _T_869 = idxHit[3] | idxHit[4]; // @[Misc.scala 182:16]
  assign _T_871 = idxHit[3] & idxHit[4]; // @[Misc.scala 182:61]
  assign _T_878 = idxHit[5] | idxHit[6]; // @[Misc.scala 182:16]
  assign _T_880 = idxHit[5] & idxHit[6]; // @[Misc.scala 182:61]
  assign _T_882 = _T_869 | _T_878; // @[Misc.scala 182:16]
  assign _T_883 = _T_871 | _T_880; // @[Misc.scala 182:37]
  assign _T_884 = _T_869 & _T_878; // @[Misc.scala 182:61]
  assign _T_885 = _T_883 | _T_884; // @[Misc.scala 182:49]
  assign _T_886 = _T_859 | _T_882; // @[Misc.scala 182:16]
  assign _T_887 = _T_862 | _T_885; // @[Misc.scala 182:37]
  assign _T_888 = _T_859 & _T_882; // @[Misc.scala 182:61]
  assign _T_889 = _T_887 | _T_888; // @[Misc.scala 182:49]
  assign _T_899 = idxHit[8] | idxHit[9]; // @[Misc.scala 182:16]
  assign _T_901 = idxHit[8] & idxHit[9]; // @[Misc.scala 182:61]
  assign _T_903 = idxHit[7] | _T_899; // @[Misc.scala 182:16]
  assign _T_905 = idxHit[7] & _T_899; // @[Misc.scala 182:61]
  assign _T_906 = _T_901 | _T_905; // @[Misc.scala 182:49]
  assign _T_913 = idxHit[10] | idxHit[11]; // @[Misc.scala 182:16]
  assign _T_915 = idxHit[10] & idxHit[11]; // @[Misc.scala 182:61]
  assign _T_922 = idxHit[12] | idxHit[13]; // @[Misc.scala 182:16]
  assign _T_924 = idxHit[12] & idxHit[13]; // @[Misc.scala 182:61]
  assign _T_926 = _T_913 | _T_922; // @[Misc.scala 182:16]
  assign _T_927 = _T_915 | _T_924; // @[Misc.scala 182:37]
  assign _T_928 = _T_913 & _T_922; // @[Misc.scala 182:61]
  assign _T_929 = _T_927 | _T_928; // @[Misc.scala 182:49]
  assign _T_930 = _T_903 | _T_926; // @[Misc.scala 182:16]
  assign _T_931 = _T_906 | _T_929; // @[Misc.scala 182:37]
  assign _T_932 = _T_903 & _T_926; // @[Misc.scala 182:61]
  assign _T_933 = _T_931 | _T_932; // @[Misc.scala 182:49]
  assign _T_934 = _T_886 | _T_930; // @[Misc.scala 182:16]
  assign _T_935 = _T_889 | _T_933; // @[Misc.scala 182:37]
  assign _T_936 = _T_886 & _T_930; // @[Misc.scala 182:61]
  assign _T_937 = _T_935 | _T_936; // @[Misc.scala 182:49]
  assign _T_948 = idxHit[15] | idxHit[16]; // @[Misc.scala 182:16]
  assign _T_950 = idxHit[15] & idxHit[16]; // @[Misc.scala 182:61]
  assign _T_952 = idxHit[14] | _T_948; // @[Misc.scala 182:16]
  assign _T_954 = idxHit[14] & _T_948; // @[Misc.scala 182:61]
  assign _T_955 = _T_950 | _T_954; // @[Misc.scala 182:49]
  assign _T_962 = idxHit[17] | idxHit[18]; // @[Misc.scala 182:16]
  assign _T_964 = idxHit[17] & idxHit[18]; // @[Misc.scala 182:61]
  assign _T_971 = idxHit[19] | idxHit[20]; // @[Misc.scala 182:16]
  assign _T_973 = idxHit[19] & idxHit[20]; // @[Misc.scala 182:61]
  assign _T_975 = _T_962 | _T_971; // @[Misc.scala 182:16]
  assign _T_976 = _T_964 | _T_973; // @[Misc.scala 182:37]
  assign _T_977 = _T_962 & _T_971; // @[Misc.scala 182:61]
  assign _T_978 = _T_976 | _T_977; // @[Misc.scala 182:49]
  assign _T_979 = _T_952 | _T_975; // @[Misc.scala 182:16]
  assign _T_980 = _T_955 | _T_978; // @[Misc.scala 182:37]
  assign _T_981 = _T_952 & _T_975; // @[Misc.scala 182:61]
  assign _T_982 = _T_980 | _T_981; // @[Misc.scala 182:49]
  assign _T_992 = idxHit[22] | idxHit[23]; // @[Misc.scala 182:16]
  assign _T_994 = idxHit[22] & idxHit[23]; // @[Misc.scala 182:61]
  assign _T_996 = idxHit[21] | _T_992; // @[Misc.scala 182:16]
  assign _T_998 = idxHit[21] & _T_992; // @[Misc.scala 182:61]
  assign _T_999 = _T_994 | _T_998; // @[Misc.scala 182:49]
  assign _T_1006 = idxHit[24] | idxHit[25]; // @[Misc.scala 182:16]
  assign _T_1008 = idxHit[24] & idxHit[25]; // @[Misc.scala 182:61]
  assign _T_1015 = idxHit[26] | idxHit[27]; // @[Misc.scala 182:16]
  assign _T_1017 = idxHit[26] & idxHit[27]; // @[Misc.scala 182:61]
  assign _T_1019 = _T_1006 | _T_1015; // @[Misc.scala 182:16]
  assign _T_1020 = _T_1008 | _T_1017; // @[Misc.scala 182:37]
  assign _T_1021 = _T_1006 & _T_1015; // @[Misc.scala 182:61]
  assign _T_1022 = _T_1020 | _T_1021; // @[Misc.scala 182:49]
  assign _T_1023 = _T_996 | _T_1019; // @[Misc.scala 182:16]
  assign _T_1024 = _T_999 | _T_1022; // @[Misc.scala 182:37]
  assign _T_1025 = _T_996 & _T_1019; // @[Misc.scala 182:61]
  assign _T_1026 = _T_1024 | _T_1025; // @[Misc.scala 182:49]
  assign _T_1027 = _T_979 | _T_1023; // @[Misc.scala 182:16]
  assign _T_1028 = _T_982 | _T_1026; // @[Misc.scala 182:37]
  assign _T_1029 = _T_979 & _T_1023; // @[Misc.scala 182:61]
  assign _T_1030 = _T_1028 | _T_1029; // @[Misc.scala 182:49]
  assign _T_1032 = _T_937 | _T_1030; // @[Misc.scala 182:37]
  assign _T_1033 = _T_934 & _T_1027; // @[Misc.scala 182:61]
  assign _T_1034 = _T_1032 | _T_1033; // @[Misc.scala 182:49]
  assign _T_1036 = isValid & ~idxHit; // @[BTB.scala 285:24]
  assign _GEN_380 = _T_1034 ? {{4'd0}, _T_1036} : _GEN_338; // @[BTB.scala 284:37]
  assign _GEN_381 = io_flush ? 32'h0 : _GEN_380; // @[BTB.scala 287:19]
  assign _T_1039 = cfiType_0 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1040 = cfiType_1 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1041 = cfiType_2 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1042 = cfiType_3 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1043 = cfiType_4 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1044 = cfiType_5 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1045 = cfiType_6 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1046 = cfiType_7 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1047 = cfiType_8 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1048 = cfiType_9 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1049 = cfiType_10 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1050 = cfiType_11 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1051 = cfiType_12 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1052 = cfiType_13 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1053 = cfiType_14 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1054 = cfiType_15 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1055 = cfiType_16 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1056 = cfiType_17 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1057 = cfiType_18 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1058 = cfiType_19 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1059 = cfiType_20 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1060 = cfiType_21 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1061 = cfiType_22 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1062 = cfiType_23 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1063 = cfiType_24 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1064 = cfiType_25 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1065 = cfiType_26 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1066 = cfiType_27 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1072 = {_T_1045,_T_1044,_T_1043,_T_1042,_T_1041,_T_1040,_T_1039}; // @[Cat.scala 29:58]
  assign _T_1079 = {_T_1052,_T_1051,_T_1050,_T_1049,_T_1048,_T_1047,_T_1046,_T_1072}; // @[Cat.scala 29:58]
  assign _T_1085 = {_T_1059,_T_1058,_T_1057,_T_1056,_T_1055,_T_1054,_T_1053}; // @[Cat.scala 29:58]
  assign _T_1093 = {_T_1066,_T_1065,_T_1064,_T_1063,_T_1062,_T_1061,_T_1060,_T_1085,_T_1079}; // @[Cat.scala 29:58]
  assign _T_1094 = idxHit & _T_1093; // @[BTB.scala 293:28]
  assign _T_1095 = |_T_1094; // @[BTB.scala 293:72]
  assign _GEN_439 = {{7'd0}, io_req_bits_addr[12:11]}; // @[BTB.scala 87:42]
  assign _T_1101 = io_req_bits_addr[10:2] ^ _GEN_439; // @[BTB.scala 87:42]
  assign _T_1102 = 8'hdd * _T_1038; // @[BTB.scala 83:12]
  assign _T_1104 = {_T_1102[7:5], 6'h0}; // @[BTB.scala 89:44]
  assign _T_1109 = {io_bht_advance_bits_bht_value,_T_1038[7:1]}; // @[Cat.scala 29:58]
  assign _GEN_440 = {{7'd0}, io_bht_update_bits_pc[12:11]}; // @[BTB.scala 87:42]
  assign _T_1114 = io_bht_update_bits_pc[10:2] ^ _GEN_440; // @[BTB.scala 87:42]
  assign _T_1115 = 8'hdd * io_bht_update_bits_prediction_history; // @[BTB.scala 83:12]
  assign _T_1117 = {_T_1115[7:5], 6'h0}; // @[BTB.scala 89:44]
  assign _T_1121 = {io_bht_update_bits_taken,io_bht_update_bits_prediction_history[7:1]}; // @[Cat.scala 29:58]
  assign _T_1096_value = _T_1037__T_1106_data; // @[BTB.scala 92:19 BTB.scala 93:15]
  assign _T_1124 = ~_T_1096_value & _T_1095; // @[BTB.scala 308:22]
  assign _T_1128 = cfiType_0 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1129 = cfiType_1 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1130 = cfiType_2 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1131 = cfiType_3 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1132 = cfiType_4 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1133 = cfiType_5 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1134 = cfiType_6 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1135 = cfiType_7 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1136 = cfiType_8 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1137 = cfiType_9 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1138 = cfiType_10 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1139 = cfiType_11 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1140 = cfiType_12 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1141 = cfiType_13 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1142 = cfiType_14 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1143 = cfiType_15 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1144 = cfiType_16 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1145 = cfiType_17 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1146 = cfiType_18 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1147 = cfiType_19 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1148 = cfiType_20 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1149 = cfiType_21 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1150 = cfiType_22 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1151 = cfiType_23 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1152 = cfiType_24 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1153 = cfiType_25 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1154 = cfiType_26 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1155 = cfiType_27 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1161 = {_T_1134,_T_1133,_T_1132,_T_1131,_T_1130,_T_1129,_T_1128}; // @[Cat.scala 29:58]
  assign _T_1168 = {_T_1141,_T_1140,_T_1139,_T_1138,_T_1137,_T_1136,_T_1135,_T_1161}; // @[Cat.scala 29:58]
  assign _T_1174 = {_T_1148,_T_1147,_T_1146,_T_1145,_T_1144,_T_1143,_T_1142}; // @[Cat.scala 29:58]
  assign _T_1182 = {_T_1155,_T_1154,_T_1153,_T_1152,_T_1151,_T_1150,_T_1149,_T_1174,_T_1168}; // @[Cat.scala 29:58]
  assign _T_1183 = idxHit & _T_1182; // @[BTB.scala 314:26]
  assign _T_1184 = |_T_1183; // @[BTB.scala 314:67]
  assign _T_1185 = _T_1125 == 3'h0; // @[BTB.scala 55:29]
  assign _GEN_399 = 3'h1 == _T_1126 ? _T_1127_1 : _T_1127_0; // @[BTB.scala 316:22]
  assign _GEN_400 = 3'h2 == _T_1126 ? _T_1127_2 : _GEN_399; // @[BTB.scala 316:22]
  assign _GEN_401 = 3'h3 == _T_1126 ? _T_1127_3 : _GEN_400; // @[BTB.scala 316:22]
  assign _GEN_402 = 3'h4 == _T_1126 ? _T_1127_4 : _GEN_401; // @[BTB.scala 316:22]
  assign _GEN_403 = 3'h5 == _T_1126 ? _T_1127_5 : _GEN_402; // @[BTB.scala 316:22]
  assign _T_1189 = ~_T_1185 & _T_1184; // @[BTB.scala 317:24]
  assign _T_1190 = io_ras_update_bits_cfiType == 2'h2; // @[BTB.scala 321:40]
  assign _T_1191 = _T_1125 < 3'h6; // @[BTB.scala 44:17]
  assign _T_1193 = _T_1125 + 3'h1; // @[BTB.scala 44:42]
  assign _T_1194 = _T_1126 < 3'h5; // @[BTB.scala 45:49]
  assign _T_1197 = _T_1126 + 3'h1; // @[BTB.scala 45:62]
  assign _T_1198 = _T_1194 ? _T_1197 : 3'h0; // @[BTB.scala 45:22]
  assign _T_1199 = io_ras_update_bits_cfiType == 2'h3; // @[BTB.scala 323:46]
  assign _T_1203 = _T_1125 - 3'h1; // @[BTB.scala 51:20]
  assign _T_1204 = _T_1126 > 3'h0; // @[BTB.scala 52:42]
  assign _T_1207 = _T_1126 - 3'h1; // @[BTB.scala 52:50]
  assign io_resp_valid = _T_477[0]; // @[BTB.scala 275:17]
  assign io_resp_bits_taken = _T_1124 ? 1'h0 : 1'h1; // @[BTB.scala 276:22 BTB.scala 308:56]
  assign io_resp_bits_bridx = _T_751 | _T_725; // @[BTB.scala 279:22]
  assign io_resp_bits_target = _T_1189 ? _GEN_403 : _T_648; // @[BTB.scala 277:23 BTB.scala 318:27]
  assign io_resp_bits_entry = {_T_651,_T_668}; // @[BTB.scala 278:22]
  assign io_resp_bits_bht_history = _T_1038; // @[BTB.scala 309:22]
  assign io_resp_bits_bht_value = _T_1037__T_1106_data; // @[BTB.scala 309:22]
  assign io_ras_head_valid = ~_T_1185; // @[BTB.scala 315:23]
  assign io_ras_head_bits = 3'h5 == _T_1126 ? _T_1127_5 : _GEN_402; // @[BTB.scala 316:22]
  assign BTB_cov_read_addr = BTB_state;
  assign BTB_cov_read_data = BTB_cov[BTB_cov_read_addr]; // @[Coverage map for BTB]
  assign BTB_cov_write_data = 1'h1;
  assign BTB_cov_write_addr = BTB_state;
  assign BTB_cov_write_mask = 1'h1;
  assign BTB_cov_write_en = 1'h1;
  assign mux_cond_0 = idxHit[20];
  assign mux_cond_1 = idxHit[3];
  assign mux_cond_2 = idxHit[26];
  assign mux_cond_3 = idxHit[4];
  assign mux_cond_4 = idxHit[27];
  assign mux_cond_5 = idxHit[12];
  assign mux_cond_6 = idxHit[5];
  assign mux_cond_7 = idxHit[24];
  assign mux_cond_8 = idxHit[21];
  assign mux_cond_9 = idxHit[9];
  assign mux_cond_10 = idxHit[17];
  assign mux_cond_11 = idxHit[8];
  assign mux_cond_12 = idxHit[0];
  assign mux_cond_13 = idxHit[25];
  assign mux_cond_14 = idxHit[10];
  assign mux_cond_15 = idxHit[2];
  assign mux_cond_16 = idxHit[7];
  assign mux_cond_17 = idxHit[18];
  assign mux_cond_18 = idxHit[14];
  assign mux_cond_19 = _T_1034;
  assign mux_cond_20 = idxHit[15];
  assign mux_cond_21 = idxHit[16];
  assign mux_cond_22 = idxHit[13];
  assign mux_cond_23 = idxHit[6];
  assign mux_cond_24 = idxHit[23];
  assign mux_cond_25 = idxHit[11];
  assign mux_cond_26 = idxHit[19];
  assign mux_cond_27 = idxHit[1];
  assign mux_cond_28 = idxHit[22];
  assign r_respPipe_bits_taken_shl = {r_respPipe_bits_taken, 6'h0};
  assign r_respPipe_bits_taken_pad = {13'h0,r_respPipe_bits_taken_shl};
  assign r_btb_updatePipe_valid_shl = {r_btb_updatePipe_valid, 16'h0};
  assign r_btb_updatePipe_valid_pad = {3'h0,r_btb_updatePipe_valid_shl};
  assign r_respPipe_valid_shl = {r_respPipe_valid, 14'h0};
  assign r_respPipe_valid_pad = {5'h0,r_respPipe_valid_shl};
  assign pageValid_shl = {pageValid, 12'h0};
  assign pageValid_pad = {2'h0,pageValid_shl};
  assign _T_1125_shl = {_T_1125, 15'h0};
  assign _T_1125_pad = {2'h0,_T_1125_shl};
  assign r_btb_updatePipe_bits_isValid_shl = {r_btb_updatePipe_bits_isValid, 10'h0};
  assign r_btb_updatePipe_bits_isValid_pad = {9'h0,r_btb_updatePipe_bits_isValid_shl};
  assign nextPageRepl_shl = {nextPageRepl, 12'h0};
  assign nextPageRepl_pad = {5'h0,nextPageRepl_shl};
  assign _T_1126_shl = {_T_1126, 16'h0};
  assign _T_1126_pad = {1'h0,_T_1126_shl};
  assign mux_cond_0_shl = {mux_cond_0, 17'h0};
  assign mux_cond_0_pad = {2'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 2'h0};
  assign mux_cond_1_pad = {17'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 3'h0};
  assign mux_cond_2_pad = {16'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 5'h0};
  assign mux_cond_3_pad = {14'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 13'h0};
  assign mux_cond_4_pad = {6'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 18'h0};
  assign mux_cond_5_pad = {1'h0,mux_cond_5_shl};
  assign mux_cond_6_shl = {mux_cond_6, 9'h0};
  assign mux_cond_6_pad = {10'h0,mux_cond_6_shl};
  assign mux_cond_7_shl = {mux_cond_7, 8'h0};
  assign mux_cond_7_pad = {11'h0,mux_cond_7_shl};
  assign mux_cond_8_shl = {mux_cond_8, 12'h0};
  assign mux_cond_8_pad = {7'h0,mux_cond_8_shl};
  assign mux_cond_9_shl = {mux_cond_9, 8'h0};
  assign mux_cond_9_pad = {11'h0,mux_cond_9_shl};
  assign mux_cond_10_shl = {mux_cond_10, 13'h0};
  assign mux_cond_10_pad = {6'h0,mux_cond_10_shl};
  assign mux_cond_11_shl = {mux_cond_11, 18'h0};
  assign mux_cond_11_pad = {1'h0,mux_cond_11_shl};
  assign mux_cond_12_shl = {mux_cond_12, 17'h0};
  assign mux_cond_12_pad = {2'h0,mux_cond_12_shl};
  assign mux_cond_13_shl = {mux_cond_13, 16'h0};
  assign mux_cond_13_pad = {3'h0,mux_cond_13_shl};
  assign mux_cond_14_shl = {mux_cond_14, 15'h0};
  assign mux_cond_14_pad = {4'h0,mux_cond_14_shl};
  assign mux_cond_15_shl = {mux_cond_15, 1'h0};
  assign mux_cond_15_pad = {18'h0,mux_cond_15_shl};
  assign mux_cond_16_shl = {mux_cond_16, 5'h0};
  assign mux_cond_16_pad = {14'h0,mux_cond_16_shl};
  assign mux_cond_17_shl = {mux_cond_17, 3'h0};
  assign mux_cond_17_pad = {16'h0,mux_cond_17_shl};
  assign mux_cond_18_shl = {mux_cond_18, 9'h0};
  assign mux_cond_18_pad = {10'h0,mux_cond_18_shl};
  assign mux_cond_19_shl = {mux_cond_19, 7'h0};
  assign mux_cond_19_pad = {12'h0,mux_cond_19_shl};
  assign mux_cond_20_shl = {mux_cond_20, 18'h0};
  assign mux_cond_20_pad = {1'h0,mux_cond_20_shl};
  assign mux_cond_21_shl = {mux_cond_21, 4'h0};
  assign mux_cond_21_pad = {15'h0,mux_cond_21_shl};
  assign mux_cond_22_shl = {mux_cond_22, 16'h0};
  assign mux_cond_22_pad = {3'h0,mux_cond_22_shl};
  assign mux_cond_23_shl = mux_cond_23;
  assign mux_cond_23_pad = {19'h0,mux_cond_23_shl};
  assign mux_cond_24_shl = {mux_cond_24, 19'h0};
  assign mux_cond_24_pad = mux_cond_24_shl;
  assign mux_cond_25_shl = {mux_cond_25, 5'h0};
  assign mux_cond_25_pad = {14'h0,mux_cond_25_shl};
  assign mux_cond_26_shl = {mux_cond_26, 15'h0};
  assign mux_cond_26_pad = {4'h0,mux_cond_26_shl};
  assign mux_cond_27_shl = {mux_cond_27, 9'h0};
  assign mux_cond_27_pad = {10'h0,mux_cond_27_shl};
  assign mux_cond_28_shl = {mux_cond_28, 12'h0};
  assign mux_cond_28_pad = {7'h0,mux_cond_28_shl};
  assign cfiType_4_shl = {cfiType_4, 12'h0};
  assign cfiType_4_pad = {6'h0,cfiType_4_shl};
  assign tgtPages_20_shl = {tgtPages_20, 7'h0};
  assign tgtPages_20_pad = {10'h0,tgtPages_20_shl};
  assign tgtPages_17_shl = {tgtPages_17, 7'h0};
  assign tgtPages_17_pad = {10'h0,tgtPages_17_shl};
  assign tgtPages_3_shl = {tgtPages_3, 7'h0};
  assign tgtPages_3_pad = {10'h0,tgtPages_3_shl};
  assign cfiType_1_shl = {cfiType_1, 12'h0};
  assign cfiType_1_pad = {6'h0,cfiType_1_shl};
  assign tgtPages_2_shl = {tgtPages_2, 7'h0};
  assign tgtPages_2_pad = {10'h0,tgtPages_2_shl};
  assign cfiType_18_shl = {cfiType_18, 12'h0};
  assign cfiType_18_pad = {6'h0,cfiType_18_shl};
  assign tgtPages_26_shl = {tgtPages_26, 7'h0};
  assign tgtPages_26_pad = {10'h0,tgtPages_26_shl};
  assign cfiType_20_shl = {cfiType_20, 12'h0};
  assign cfiType_20_pad = {6'h0,cfiType_20_shl};
  assign cfiType_22_shl = {cfiType_22, 12'h0};
  assign cfiType_22_pad = {6'h0,cfiType_22_shl};
  assign cfiType_23_shl = {cfiType_23, 12'h0};
  assign cfiType_23_pad = {6'h0,cfiType_23_shl};
  assign cfiType_0_shl = {cfiType_0, 12'h0};
  assign cfiType_0_pad = {6'h0,cfiType_0_shl};
  assign tgtPages_11_shl = {tgtPages_11, 7'h0};
  assign tgtPages_11_pad = {10'h0,tgtPages_11_shl};
  assign cfiType_7_shl = {cfiType_7, 12'h0};
  assign cfiType_7_pad = {6'h0,cfiType_7_shl};
  assign cfiType_19_shl = {cfiType_19, 12'h0};
  assign cfiType_19_pad = {6'h0,cfiType_19_shl};
  assign cfiType_17_shl = {cfiType_17, 12'h0};
  assign cfiType_17_pad = {6'h0,cfiType_17_shl};
  assign cfiType_25_shl = {cfiType_25, 12'h0};
  assign cfiType_25_pad = {6'h0,cfiType_25_shl};
  assign cfiType_3_shl = {cfiType_3, 12'h0};
  assign cfiType_3_pad = {6'h0,cfiType_3_shl};
  assign cfiType_10_shl = {cfiType_10, 12'h0};
  assign cfiType_10_pad = {6'h0,cfiType_10_shl};
  assign tgtPages_14_shl = {tgtPages_14, 7'h0};
  assign tgtPages_14_pad = {10'h0,tgtPages_14_shl};
  assign cfiType_2_shl = {cfiType_2, 12'h0};
  assign cfiType_2_pad = {6'h0,cfiType_2_shl};
  assign cfiType_16_shl = {cfiType_16, 12'h0};
  assign cfiType_16_pad = {6'h0,cfiType_16_shl};
  assign tgtPages_0_shl = {tgtPages_0, 7'h0};
  assign tgtPages_0_pad = {10'h0,tgtPages_0_shl};
  assign tgtPages_21_shl = {tgtPages_21, 7'h0};
  assign tgtPages_21_pad = {10'h0,tgtPages_21_shl};
  assign tgtPages_5_shl = {tgtPages_5, 7'h0};
  assign tgtPages_5_pad = {10'h0,tgtPages_5_shl};
  assign tgtPages_4_shl = {tgtPages_4, 7'h0};
  assign tgtPages_4_pad = {10'h0,tgtPages_4_shl};
  assign cfiType_9_shl = {cfiType_9, 12'h0};
  assign cfiType_9_pad = {6'h0,cfiType_9_shl};
  assign tgtPages_25_shl = {tgtPages_25, 7'h0};
  assign tgtPages_25_pad = {10'h0,tgtPages_25_shl};
  assign cfiType_8_shl = {cfiType_8, 12'h0};
  assign cfiType_8_pad = {6'h0,cfiType_8_shl};
  assign tgtPages_24_shl = {tgtPages_24, 7'h0};
  assign tgtPages_24_pad = {10'h0,tgtPages_24_shl};
  assign cfiType_26_shl = {cfiType_26, 12'h0};
  assign cfiType_26_pad = {6'h0,cfiType_26_shl};
  assign tgtPages_13_shl = {tgtPages_13, 7'h0};
  assign tgtPages_13_pad = {10'h0,tgtPages_13_shl};
  assign cfiType_14_shl = {cfiType_14, 12'h0};
  assign cfiType_14_pad = {6'h0,cfiType_14_shl};
  assign cfiType_11_shl = {cfiType_11, 12'h0};
  assign cfiType_11_pad = {6'h0,cfiType_11_shl};
  assign tgtPages_16_shl = {tgtPages_16, 7'h0};
  assign tgtPages_16_pad = {10'h0,tgtPages_16_shl};
  assign cfiType_15_shl = {cfiType_15, 12'h0};
  assign cfiType_15_pad = {6'h0,cfiType_15_shl};
  assign cfiType_24_shl = {cfiType_24, 12'h0};
  assign cfiType_24_pad = {6'h0,cfiType_24_shl};
  assign tgtPages_18_shl = {tgtPages_18, 7'h0};
  assign tgtPages_18_pad = {10'h0,tgtPages_18_shl};
  assign cfiType_21_shl = {cfiType_21, 12'h0};
  assign cfiType_21_pad = {6'h0,cfiType_21_shl};
  assign tgtPages_12_shl = {tgtPages_12, 7'h0};
  assign tgtPages_12_pad = {10'h0,tgtPages_12_shl};
  assign tgtPages_10_shl = {tgtPages_10, 7'h0};
  assign tgtPages_10_pad = {10'h0,tgtPages_10_shl};
  assign tgtPages_15_shl = {tgtPages_15, 7'h0};
  assign tgtPages_15_pad = {10'h0,tgtPages_15_shl};
  assign tgtPages_22_shl = {tgtPages_22, 7'h0};
  assign tgtPages_22_pad = {10'h0,tgtPages_22_shl};
  assign tgtPages_19_shl = {tgtPages_19, 7'h0};
  assign tgtPages_19_pad = {10'h0,tgtPages_19_shl};
  assign cfiType_13_shl = {cfiType_13, 12'h0};
  assign cfiType_13_pad = {6'h0,cfiType_13_shl};
  assign cfiType_6_shl = {cfiType_6, 12'h0};
  assign cfiType_6_pad = {6'h0,cfiType_6_shl};
  assign tgtPages_6_shl = {tgtPages_6, 7'h0};
  assign tgtPages_6_pad = {10'h0,tgtPages_6_shl};
  assign cfiType_27_shl = {cfiType_27, 12'h0};
  assign cfiType_27_pad = {6'h0,cfiType_27_shl};
  assign tgtPages_23_shl = {tgtPages_23, 7'h0};
  assign tgtPages_23_pad = {10'h0,tgtPages_23_shl};
  assign cfiType_12_shl = {cfiType_12, 12'h0};
  assign cfiType_12_pad = {6'h0,cfiType_12_shl};
  assign tgtPages_8_shl = {tgtPages_8, 7'h0};
  assign tgtPages_8_pad = {10'h0,tgtPages_8_shl};
  assign tgtPages_1_shl = {tgtPages_1, 7'h0};
  assign tgtPages_1_pad = {10'h0,tgtPages_1_shl};
  assign tgtPages_9_shl = {tgtPages_9, 7'h0};
  assign tgtPages_9_pad = {10'h0,tgtPages_9_shl};
  assign cfiType_5_shl = {cfiType_5, 12'h0};
  assign cfiType_5_pad = {6'h0,cfiType_5_shl};
  assign tgtPages_7_shl = {tgtPages_7, 7'h0};
  assign tgtPages_7_pad = {10'h0,tgtPages_7_shl};
  assign tgtPages_27_shl = {tgtPages_27, 7'h0};
  assign tgtPages_27_pad = {10'h0,tgtPages_27_shl};
  assign BTB_xor31 = r_respPipe_bits_taken_pad ^ r_btb_updatePipe_valid_pad;
  assign BTB_xor66 = pageValid_pad ^ _T_1125_pad;
  assign BTB_xor32 = r_respPipe_valid_pad ^ BTB_xor66;
  assign BTB_xor15 = BTB_xor31 ^ BTB_xor32;
  assign BTB_xor68 = nextPageRepl_pad ^ _T_1126_pad;
  assign BTB_xor33 = r_btb_updatePipe_bits_isValid_pad ^ BTB_xor68;
  assign BTB_xor70 = mux_cond_1_pad ^ mux_cond_2_pad;
  assign BTB_xor34 = mux_cond_0_pad ^ BTB_xor70;
  assign BTB_xor16 = BTB_xor33 ^ BTB_xor34;
  assign BTB_xor7 = BTB_xor15 ^ BTB_xor16;
  assign BTB_xor72 = mux_cond_4_pad ^ mux_cond_5_pad;
  assign BTB_xor35 = mux_cond_3_pad ^ BTB_xor72;
  assign BTB_xor74 = mux_cond_7_pad ^ mux_cond_8_pad;
  assign BTB_xor36 = mux_cond_6_pad ^ BTB_xor74;
  assign BTB_xor17 = BTB_xor35 ^ BTB_xor36;
  assign BTB_xor76 = mux_cond_10_pad ^ mux_cond_11_pad;
  assign BTB_xor37 = mux_cond_9_pad ^ BTB_xor76;
  assign BTB_xor78 = mux_cond_13_pad ^ mux_cond_14_pad;
  assign BTB_xor38 = mux_cond_12_pad ^ BTB_xor78;
  assign BTB_xor18 = BTB_xor37 ^ BTB_xor38;
  assign BTB_xor8 = BTB_xor17 ^ BTB_xor18;
  assign BTB_xor3 = BTB_xor7 ^ BTB_xor8;
  assign BTB_xor39 = mux_cond_15_pad ^ mux_cond_16_pad;
  assign BTB_xor82 = mux_cond_18_pad ^ mux_cond_19_pad;
  assign BTB_xor40 = mux_cond_17_pad ^ BTB_xor82;
  assign BTB_xor19 = BTB_xor39 ^ BTB_xor40;
  assign BTB_xor84 = mux_cond_21_pad ^ mux_cond_22_pad;
  assign BTB_xor41 = mux_cond_20_pad ^ BTB_xor84;
  assign BTB_xor86 = mux_cond_24_pad ^ mux_cond_25_pad;
  assign BTB_xor42 = mux_cond_23_pad ^ BTB_xor86;
  assign BTB_xor20 = BTB_xor41 ^ BTB_xor42;
  assign BTB_xor9 = BTB_xor19 ^ BTB_xor20;
  assign BTB_xor88 = mux_cond_27_pad ^ mux_cond_28_pad;
  assign BTB_xor43 = mux_cond_26_pad ^ BTB_xor88;
  assign BTB_xor90 = tgtPages_20_pad ^ tgtPages_17_pad;
  assign BTB_xor44 = cfiType_4_pad ^ BTB_xor90;
  assign BTB_xor21 = BTB_xor43 ^ BTB_xor44;
  assign BTB_xor92 = cfiType_1_pad ^ tgtPages_2_pad;
  assign BTB_xor45 = tgtPages_3_pad ^ BTB_xor92;
  assign BTB_xor94 = tgtPages_26_pad ^ cfiType_20_pad;
  assign BTB_xor46 = cfiType_18_pad ^ BTB_xor94;
  assign BTB_xor22 = BTB_xor45 ^ BTB_xor46;
  assign BTB_xor10 = BTB_xor21 ^ BTB_xor22;
  assign BTB_xor4 = BTB_xor9 ^ BTB_xor10;
  assign BTB_xor1 = BTB_xor3 ^ BTB_xor4;
  assign BTB_xor47 = cfiType_22_pad ^ cfiType_23_pad;
  assign BTB_xor98 = tgtPages_11_pad ^ cfiType_7_pad;
  assign BTB_xor48 = cfiType_0_pad ^ BTB_xor98;
  assign BTB_xor23 = BTB_xor47 ^ BTB_xor48;
  assign BTB_xor100 = cfiType_17_pad ^ cfiType_25_pad;
  assign BTB_xor49 = cfiType_19_pad ^ BTB_xor100;
  assign BTB_xor102 = cfiType_10_pad ^ tgtPages_14_pad;
  assign BTB_xor50 = cfiType_3_pad ^ BTB_xor102;
  assign BTB_xor24 = BTB_xor49 ^ BTB_xor50;
  assign BTB_xor11 = BTB_xor23 ^ BTB_xor24;
  assign BTB_xor104 = cfiType_16_pad ^ tgtPages_0_pad;
  assign BTB_xor51 = cfiType_2_pad ^ BTB_xor104;
  assign BTB_xor106 = tgtPages_5_pad ^ tgtPages_4_pad;
  assign BTB_xor52 = tgtPages_21_pad ^ BTB_xor106;
  assign BTB_xor25 = BTB_xor51 ^ BTB_xor52;
  assign BTB_xor108 = tgtPages_25_pad ^ cfiType_8_pad;
  assign BTB_xor53 = cfiType_9_pad ^ BTB_xor108;
  assign BTB_xor110 = cfiType_26_pad ^ tgtPages_13_pad;
  assign BTB_xor54 = tgtPages_24_pad ^ BTB_xor110;
  assign BTB_xor26 = BTB_xor53 ^ BTB_xor54;
  assign BTB_xor12 = BTB_xor25 ^ BTB_xor26;
  assign BTB_xor5 = BTB_xor11 ^ BTB_xor12;
  assign BTB_xor112 = cfiType_11_pad ^ tgtPages_16_pad;
  assign BTB_xor55 = cfiType_14_pad ^ BTB_xor112;
  assign BTB_xor114 = cfiType_24_pad ^ tgtPages_18_pad;
  assign BTB_xor56 = cfiType_15_pad ^ BTB_xor114;
  assign BTB_xor27 = BTB_xor55 ^ BTB_xor56;
  assign BTB_xor116 = tgtPages_12_pad ^ tgtPages_10_pad;
  assign BTB_xor57 = cfiType_21_pad ^ BTB_xor116;
  assign BTB_xor118 = tgtPages_22_pad ^ tgtPages_19_pad;
  assign BTB_xor58 = tgtPages_15_pad ^ BTB_xor118;
  assign BTB_xor28 = BTB_xor57 ^ BTB_xor58;
  assign BTB_xor13 = BTB_xor27 ^ BTB_xor28;
  assign BTB_xor120 = cfiType_6_pad ^ tgtPages_6_pad;
  assign BTB_xor59 = cfiType_13_pad ^ BTB_xor120;
  assign BTB_xor122 = tgtPages_23_pad ^ cfiType_12_pad;
  assign BTB_xor60 = cfiType_27_pad ^ BTB_xor122;
  assign BTB_xor29 = BTB_xor59 ^ BTB_xor60;
  assign BTB_xor124 = tgtPages_1_pad ^ tgtPages_9_pad;
  assign BTB_xor61 = tgtPages_8_pad ^ BTB_xor124;
  assign BTB_xor126 = tgtPages_7_pad ^ tgtPages_27_pad;
  assign BTB_xor62 = cfiType_5_pad ^ BTB_xor126;
  assign BTB_xor30 = BTB_xor61 ^ BTB_xor62;
  assign BTB_xor14 = BTB_xor29 ^ BTB_xor30;
  assign BTB_xor6 = BTB_xor13 ^ BTB_xor14;
  assign BTB_xor2 = BTB_xor5 ^ BTB_xor6;
  assign BTB_xor0 = BTB_xor1 ^ BTB_xor2;
  assign io_covSum = BTB_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    _T_1037[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  idxs_0 = _RAND_1[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  idxs_1 = _RAND_2[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  idxs_2 = _RAND_3[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  idxs_3 = _RAND_4[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  idxs_4 = _RAND_5[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  idxs_5 = _RAND_6[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  idxs_6 = _RAND_7[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  idxs_7 = _RAND_8[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idxs_8 = _RAND_9[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idxs_9 = _RAND_10[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  idxs_10 = _RAND_11[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  idxs_11 = _RAND_12[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  idxs_12 = _RAND_13[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  idxs_13 = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  idxs_14 = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  idxs_15 = _RAND_16[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  idxs_16 = _RAND_17[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  idxs_17 = _RAND_18[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  idxs_18 = _RAND_19[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  idxs_19 = _RAND_20[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  idxs_20 = _RAND_21[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  idxs_21 = _RAND_22[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  idxs_22 = _RAND_23[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  idxs_23 = _RAND_24[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  idxs_24 = _RAND_25[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  idxs_25 = _RAND_26[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  idxs_26 = _RAND_27[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  idxs_27 = _RAND_28[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  idxPages_0 = _RAND_29[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  idxPages_1 = _RAND_30[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  idxPages_2 = _RAND_31[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  idxPages_3 = _RAND_32[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  idxPages_4 = _RAND_33[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  idxPages_5 = _RAND_34[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  idxPages_6 = _RAND_35[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  idxPages_7 = _RAND_36[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  idxPages_8 = _RAND_37[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  idxPages_9 = _RAND_38[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  idxPages_10 = _RAND_39[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  idxPages_11 = _RAND_40[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  idxPages_12 = _RAND_41[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  idxPages_13 = _RAND_42[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  idxPages_14 = _RAND_43[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  idxPages_15 = _RAND_44[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  idxPages_16 = _RAND_45[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  idxPages_17 = _RAND_46[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  idxPages_18 = _RAND_47[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  idxPages_19 = _RAND_48[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  idxPages_20 = _RAND_49[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  idxPages_21 = _RAND_50[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  idxPages_22 = _RAND_51[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  idxPages_23 = _RAND_52[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  idxPages_24 = _RAND_53[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  idxPages_25 = _RAND_54[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  idxPages_26 = _RAND_55[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  idxPages_27 = _RAND_56[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  tgts_0 = _RAND_57[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  tgts_1 = _RAND_58[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  tgts_2 = _RAND_59[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  tgts_3 = _RAND_60[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  tgts_4 = _RAND_61[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  tgts_5 = _RAND_62[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  tgts_6 = _RAND_63[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  tgts_7 = _RAND_64[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  tgts_8 = _RAND_65[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  tgts_9 = _RAND_66[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  tgts_10 = _RAND_67[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  tgts_11 = _RAND_68[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  tgts_12 = _RAND_69[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  tgts_13 = _RAND_70[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  tgts_14 = _RAND_71[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  tgts_15 = _RAND_72[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  tgts_16 = _RAND_73[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  tgts_17 = _RAND_74[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  tgts_18 = _RAND_75[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  tgts_19 = _RAND_76[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  tgts_20 = _RAND_77[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  tgts_21 = _RAND_78[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  tgts_22 = _RAND_79[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  tgts_23 = _RAND_80[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  tgts_24 = _RAND_81[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  tgts_25 = _RAND_82[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  tgts_26 = _RAND_83[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  tgts_27 = _RAND_84[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  tgtPages_0 = _RAND_85[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  tgtPages_1 = _RAND_86[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  tgtPages_2 = _RAND_87[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  tgtPages_3 = _RAND_88[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  tgtPages_4 = _RAND_89[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  tgtPages_5 = _RAND_90[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  tgtPages_6 = _RAND_91[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  tgtPages_7 = _RAND_92[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  tgtPages_8 = _RAND_93[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  tgtPages_9 = _RAND_94[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  tgtPages_10 = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  tgtPages_11 = _RAND_96[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  tgtPages_12 = _RAND_97[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  tgtPages_13 = _RAND_98[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  tgtPages_14 = _RAND_99[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  tgtPages_15 = _RAND_100[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  tgtPages_16 = _RAND_101[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  tgtPages_17 = _RAND_102[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  tgtPages_18 = _RAND_103[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  tgtPages_19 = _RAND_104[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  tgtPages_20 = _RAND_105[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  tgtPages_21 = _RAND_106[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  tgtPages_22 = _RAND_107[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  tgtPages_23 = _RAND_108[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  tgtPages_24 = _RAND_109[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  tgtPages_25 = _RAND_110[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  tgtPages_26 = _RAND_111[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  tgtPages_27 = _RAND_112[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  pages_0 = _RAND_113[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  pages_1 = _RAND_114[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  pages_2 = _RAND_115[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  pages_3 = _RAND_116[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  pages_4 = _RAND_117[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  pages_5 = _RAND_118[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  pageValid = _RAND_119[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  isValid = _RAND_120[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  cfiType_0 = _RAND_121[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  cfiType_1 = _RAND_122[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  cfiType_2 = _RAND_123[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  cfiType_3 = _RAND_124[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  cfiType_4 = _RAND_125[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  cfiType_5 = _RAND_126[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  cfiType_6 = _RAND_127[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  cfiType_7 = _RAND_128[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  cfiType_8 = _RAND_129[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  cfiType_9 = _RAND_130[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  cfiType_10 = _RAND_131[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  cfiType_11 = _RAND_132[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  cfiType_12 = _RAND_133[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  cfiType_13 = _RAND_134[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  cfiType_14 = _RAND_135[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  cfiType_15 = _RAND_136[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  cfiType_16 = _RAND_137[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  cfiType_17 = _RAND_138[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  cfiType_18 = _RAND_139[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  cfiType_19 = _RAND_140[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  cfiType_20 = _RAND_141[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  cfiType_21 = _RAND_142[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  cfiType_22 = _RAND_143[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  cfiType_23 = _RAND_144[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  cfiType_24 = _RAND_145[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  cfiType_25 = _RAND_146[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  cfiType_26 = _RAND_147[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  cfiType_27 = _RAND_148[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  brIdx_0 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  brIdx_1 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  brIdx_2 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  brIdx_3 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  brIdx_4 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  brIdx_5 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  brIdx_6 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  brIdx_7 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  brIdx_8 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  brIdx_9 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  brIdx_10 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  brIdx_11 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  brIdx_12 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  brIdx_13 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  brIdx_14 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  brIdx_15 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  brIdx_16 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  brIdx_17 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  brIdx_18 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  brIdx_19 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  brIdx_20 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  brIdx_21 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  brIdx_22 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  brIdx_23 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  brIdx_24 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  brIdx_25 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  brIdx_26 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  brIdx_27 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  r_btb_updatePipe_valid = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  r_btb_updatePipe_bits_prediction_entry = _RAND_178[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {2{`RANDOM}};
  r_btb_updatePipe_bits_pc = _RAND_179[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  r_btb_updatePipe_bits_isValid = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {2{`RANDOM}};
  r_btb_updatePipe_bits_br_pc = _RAND_181[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  r_btb_updatePipe_bits_cfiType = _RAND_182[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  nextPageRepl = _RAND_183[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_123 = _RAND_184[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  r_respPipe_valid = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  r_respPipe_bits_taken = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  r_respPipe_bits_entry = _RAND_187[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_1038 = _RAND_188[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_1125 = _RAND_189[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_1126 = _RAND_190[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {2{`RANDOM}};
  _T_1127_0 = _RAND_191[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {2{`RANDOM}};
  _T_1127_1 = _RAND_192[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {2{`RANDOM}};
  _T_1127_2 = _RAND_193[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {2{`RANDOM}};
  _T_1127_3 = _RAND_194[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {2{`RANDOM}};
  _T_1127_4 = _RAND_195[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {2{`RANDOM}};
  _T_1127_5 = _RAND_196[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  BTB_state = _RAND_197[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    BTB_cov[initvar] = _RAND_198[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  BTB_covSum = _RAND_199[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_1037__T_1119_en & _T_1037__T_1119_mask) begin
      _T_1037[_T_1037__T_1119_addr] <= _T_1037__T_1119_data; // @[BTB.scala 113:26]
    end
    if (metaReset) begin
      idxs_0 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h0 == waddr) begin
        idxs_0 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_1 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1 == waddr) begin
        idxs_1 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_2 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h2 == waddr) begin
        idxs_2 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_3 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h3 == waddr) begin
        idxs_3 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_4 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h4 == waddr) begin
        idxs_4 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_5 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h5 == waddr) begin
        idxs_5 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_6 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h6 == waddr) begin
        idxs_6 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_7 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h7 == waddr) begin
        idxs_7 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_8 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h8 == waddr) begin
        idxs_8 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_9 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h9 == waddr) begin
        idxs_9 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_10 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'ha == waddr) begin
        idxs_10 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_11 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hb == waddr) begin
        idxs_11 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_12 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hc == waddr) begin
        idxs_12 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_13 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hd == waddr) begin
        idxs_13 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_14 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'he == waddr) begin
        idxs_14 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_15 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hf == waddr) begin
        idxs_15 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_16 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h10 == waddr) begin
        idxs_16 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_17 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h11 == waddr) begin
        idxs_17 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_18 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h12 == waddr) begin
        idxs_18 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_19 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h13 == waddr) begin
        idxs_19 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_20 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h14 == waddr) begin
        idxs_20 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_21 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h15 == waddr) begin
        idxs_21 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_22 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h16 == waddr) begin
        idxs_22 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_23 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h17 == waddr) begin
        idxs_23 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_24 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h18 == waddr) begin
        idxs_24 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_25 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h19 == waddr) begin
        idxs_25 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_26 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1a == waddr) begin
        idxs_26 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_27 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1b == waddr) begin
        idxs_27 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxPages_0 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h0 == waddr) begin
        idxPages_0 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_1 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1 == waddr) begin
        idxPages_1 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_2 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h2 == waddr) begin
        idxPages_2 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_3 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h3 == waddr) begin
        idxPages_3 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_4 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h4 == waddr) begin
        idxPages_4 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_5 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h5 == waddr) begin
        idxPages_5 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_6 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h6 == waddr) begin
        idxPages_6 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_7 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h7 == waddr) begin
        idxPages_7 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_8 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h8 == waddr) begin
        idxPages_8 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_9 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h9 == waddr) begin
        idxPages_9 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_10 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'ha == waddr) begin
        idxPages_10 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_11 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hb == waddr) begin
        idxPages_11 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_12 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hc == waddr) begin
        idxPages_12 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_13 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hd == waddr) begin
        idxPages_13 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_14 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'he == waddr) begin
        idxPages_14 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_15 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hf == waddr) begin
        idxPages_15 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_16 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h10 == waddr) begin
        idxPages_16 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_17 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h11 == waddr) begin
        idxPages_17 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_18 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h12 == waddr) begin
        idxPages_18 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_19 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h13 == waddr) begin
        idxPages_19 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_20 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h14 == waddr) begin
        idxPages_20 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_21 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h15 == waddr) begin
        idxPages_21 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_22 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h16 == waddr) begin
        idxPages_22 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_23 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h17 == waddr) begin
        idxPages_23 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_24 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h18 == waddr) begin
        idxPages_24 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_25 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h19 == waddr) begin
        idxPages_25 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_26 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1a == waddr) begin
        idxPages_26 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      idxPages_27 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1b == waddr) begin
        idxPages_27 <= _T_368[2:0];
      end
    end
    if (metaReset) begin
      tgts_0 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h0 == waddr) begin
        tgts_0 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_1 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1 == waddr) begin
        tgts_1 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_2 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h2 == waddr) begin
        tgts_2 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_3 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h3 == waddr) begin
        tgts_3 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_4 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h4 == waddr) begin
        tgts_4 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_5 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h5 == waddr) begin
        tgts_5 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_6 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h6 == waddr) begin
        tgts_6 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_7 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h7 == waddr) begin
        tgts_7 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_8 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h8 == waddr) begin
        tgts_8 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_9 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h9 == waddr) begin
        tgts_9 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_10 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'ha == waddr) begin
        tgts_10 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_11 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hb == waddr) begin
        tgts_11 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_12 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hc == waddr) begin
        tgts_12 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_13 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hd == waddr) begin
        tgts_13 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_14 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'he == waddr) begin
        tgts_14 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_15 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hf == waddr) begin
        tgts_15 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_16 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h10 == waddr) begin
        tgts_16 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_17 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h11 == waddr) begin
        tgts_17 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_18 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h12 == waddr) begin
        tgts_18 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_19 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h13 == waddr) begin
        tgts_19 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_20 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h14 == waddr) begin
        tgts_20 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_21 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h15 == waddr) begin
        tgts_21 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_22 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h16 == waddr) begin
        tgts_22 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_23 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h17 == waddr) begin
        tgts_23 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_24 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h18 == waddr) begin
        tgts_24 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_25 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h19 == waddr) begin
        tgts_25 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_26 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1a == waddr) begin
        tgts_26 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_27 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1b == waddr) begin
        tgts_27 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgtPages_0 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h0 == waddr) begin
        tgtPages_0 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_1 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1 == waddr) begin
        tgtPages_1 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_2 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h2 == waddr) begin
        tgtPages_2 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_3 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h3 == waddr) begin
        tgtPages_3 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_4 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h4 == waddr) begin
        tgtPages_4 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_5 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h5 == waddr) begin
        tgtPages_5 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_6 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h6 == waddr) begin
        tgtPages_6 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_7 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h7 == waddr) begin
        tgtPages_7 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_8 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h8 == waddr) begin
        tgtPages_8 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_9 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h9 == waddr) begin
        tgtPages_9 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_10 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'ha == waddr) begin
        tgtPages_10 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_11 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hb == waddr) begin
        tgtPages_11 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_12 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hc == waddr) begin
        tgtPages_12 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_13 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hd == waddr) begin
        tgtPages_13 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_14 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'he == waddr) begin
        tgtPages_14 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_15 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hf == waddr) begin
        tgtPages_15 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_16 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h10 == waddr) begin
        tgtPages_16 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_17 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h11 == waddr) begin
        tgtPages_17 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_18 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h12 == waddr) begin
        tgtPages_18 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_19 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h13 == waddr) begin
        tgtPages_19 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_20 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h14 == waddr) begin
        tgtPages_20 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_21 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h15 == waddr) begin
        tgtPages_21 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_22 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h16 == waddr) begin
        tgtPages_22 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_23 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h17 == waddr) begin
        tgtPages_23 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_24 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h18 == waddr) begin
        tgtPages_24 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_25 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h19 == waddr) begin
        tgtPages_25 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_26 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1a == waddr) begin
        tgtPages_26 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_27 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1b == waddr) begin
        tgtPages_27 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      pages_0 <= 25'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (_T_376[0]) begin
        if (~idxPageUpdate[0]) begin
          pages_0 <= r_btb_updatePipe_bits_pc[38:14];
        end else begin
          pages_0 <= io_req_bits_addr[38:14];
        end
      end
    end
    if (metaReset) begin
      pages_1 <= 25'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (_T_383[1]) begin
        if (~idxPageUpdate[0]) begin
          pages_1 <= io_req_bits_addr[38:14];
        end else begin
          pages_1 <= r_btb_updatePipe_bits_pc[38:14];
        end
      end
    end
    if (metaReset) begin
      pages_2 <= 25'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (_T_376[2]) begin
        if (~idxPageUpdate[0]) begin
          pages_2 <= r_btb_updatePipe_bits_pc[38:14];
        end else begin
          pages_2 <= io_req_bits_addr[38:14];
        end
      end
    end
    if (metaReset) begin
      pages_3 <= 25'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (_T_383[3]) begin
        if (~idxPageUpdate[0]) begin
          pages_3 <= io_req_bits_addr[38:14];
        end else begin
          pages_3 <= r_btb_updatePipe_bits_pc[38:14];
        end
      end
    end
    if (metaReset) begin
      pages_4 <= 25'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (_T_376[4]) begin
        if (~idxPageUpdate[0]) begin
          pages_4 <= r_btb_updatePipe_bits_pc[38:14];
        end else begin
          pages_4 <= io_req_bits_addr[38:14];
        end
      end
    end
    if (metaReset) begin
      pages_5 <= 25'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (_T_383[5]) begin
        if (~idxPageUpdate[0]) begin
          pages_5 <= io_req_bits_addr[38:14];
        end else begin
          pages_5 <= r_btb_updatePipe_bits_pc[38:14];
        end
      end
    end
    if (metaReset) begin
      pageValid <= 6'h0;
    end else if (reset) begin
      pageValid <= 6'h0;
    end else begin
      pageValid <= _GEN_373[5:0];
    end
    if (metaReset) begin
      isValid <= 28'h0;
    end else if (reset) begin
      isValid <= 28'h0;
    end else begin
      isValid <= _GEN_381[27:0];
    end
    if (metaReset) begin
      cfiType_0 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h0 == waddr) begin
        cfiType_0 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_1 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1 == waddr) begin
        cfiType_1 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_2 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h2 == waddr) begin
        cfiType_2 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_3 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h3 == waddr) begin
        cfiType_3 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_4 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h4 == waddr) begin
        cfiType_4 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_5 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h5 == waddr) begin
        cfiType_5 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_6 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h6 == waddr) begin
        cfiType_6 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_7 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h7 == waddr) begin
        cfiType_7 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_8 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h8 == waddr) begin
        cfiType_8 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_9 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h9 == waddr) begin
        cfiType_9 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_10 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'ha == waddr) begin
        cfiType_10 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_11 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hb == waddr) begin
        cfiType_11 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_12 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hc == waddr) begin
        cfiType_12 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_13 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hd == waddr) begin
        cfiType_13 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_14 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'he == waddr) begin
        cfiType_14 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_15 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hf == waddr) begin
        cfiType_15 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_16 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h10 == waddr) begin
        cfiType_16 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_17 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h11 == waddr) begin
        cfiType_17 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_18 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h12 == waddr) begin
        cfiType_18 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_19 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h13 == waddr) begin
        cfiType_19 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_20 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h14 == waddr) begin
        cfiType_20 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_21 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h15 == waddr) begin
        cfiType_21 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_22 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h16 == waddr) begin
        cfiType_22 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_23 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h17 == waddr) begin
        cfiType_23 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_24 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h18 == waddr) begin
        cfiType_24 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_25 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h19 == waddr) begin
        cfiType_25 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_26 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1a == waddr) begin
        cfiType_26 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_27 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1b == waddr) begin
        cfiType_27 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      brIdx_0 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h0 == waddr) begin
        brIdx_0 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_1 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1 == waddr) begin
        brIdx_1 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_2 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h2 == waddr) begin
        brIdx_2 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_3 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h3 == waddr) begin
        brIdx_3 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_4 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h4 == waddr) begin
        brIdx_4 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_5 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h5 == waddr) begin
        brIdx_5 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_6 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h6 == waddr) begin
        brIdx_6 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_7 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h7 == waddr) begin
        brIdx_7 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_8 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h8 == waddr) begin
        brIdx_8 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_9 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h9 == waddr) begin
        brIdx_9 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_10 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'ha == waddr) begin
        brIdx_10 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_11 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hb == waddr) begin
        brIdx_11 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_12 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hc == waddr) begin
        brIdx_12 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_13 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hd == waddr) begin
        brIdx_13 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_14 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'he == waddr) begin
        brIdx_14 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_15 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hf == waddr) begin
        brIdx_15 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_16 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h10 == waddr) begin
        brIdx_16 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_17 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h11 == waddr) begin
        brIdx_17 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_18 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h12 == waddr) begin
        brIdx_18 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_19 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h13 == waddr) begin
        brIdx_19 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_20 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h14 == waddr) begin
        brIdx_20 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_21 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h15 == waddr) begin
        brIdx_21 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_22 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h16 == waddr) begin
        brIdx_22 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_23 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h17 == waddr) begin
        brIdx_23 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_24 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h18 == waddr) begin
        brIdx_24 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_25 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h19 == waddr) begin
        brIdx_25 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_26 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1a == waddr) begin
        brIdx_26 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_27 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1b == waddr) begin
        brIdx_27 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      r_btb_updatePipe_valid <= 1'h0;
    end else if (reset) begin
      r_btb_updatePipe_valid <= 1'h0;
    end else begin
      r_btb_updatePipe_valid <= io_btb_update_valid;
    end
    if (metaReset) begin
      r_btb_updatePipe_bits_prediction_entry <= 5'h0;
    end else if (io_btb_update_valid) begin
      r_btb_updatePipe_bits_prediction_entry <= io_btb_update_bits_prediction_entry;
    end
    if (metaReset) begin
      r_btb_updatePipe_bits_pc <= 39'h0;
    end else if (io_btb_update_valid) begin
      r_btb_updatePipe_bits_pc <= io_btb_update_bits_pc;
    end
    if (metaReset) begin
      r_btb_updatePipe_bits_isValid <= 1'h0;
    end else if (io_btb_update_valid) begin
      r_btb_updatePipe_bits_isValid <= io_btb_update_bits_isValid;
    end
    if (metaReset) begin
      r_btb_updatePipe_bits_br_pc <= 39'h0;
    end else if (io_btb_update_valid) begin
      r_btb_updatePipe_bits_br_pc <= io_btb_update_bits_br_pc;
    end
    if (metaReset) begin
      r_btb_updatePipe_bits_cfiType <= 2'h0;
    end else if (io_btb_update_valid) begin
      r_btb_updatePipe_bits_cfiType <= io_btb_update_bits_cfiType;
    end
    if (metaReset) begin
      nextPageRepl <= 3'h0;
    end else if (_T_115) begin
      if (_T_120) begin
        nextPageRepl <= {{2'd0}, _T_119[0]};
      end else begin
        nextPageRepl <= _T_119;
      end
    end
    if (metaReset) begin
      _T_123 <= 27'h0;
    end else if (_T_204) begin
      _T_123 <= _T_364;
    end
    if (metaReset) begin
      r_respPipe_valid <= 1'h0;
    end else if (reset) begin
      r_respPipe_valid <= 1'h0;
    end else begin
      r_respPipe_valid <= io_resp_valid;
    end
    if (metaReset) begin
      r_respPipe_bits_taken <= 1'h0;
    end else if (io_resp_valid) begin
      r_respPipe_bits_taken <= io_resp_bits_taken;
    end
    if (metaReset) begin
      r_respPipe_bits_entry <= 5'h0;
    end else if (io_resp_valid) begin
      r_respPipe_bits_entry <= io_resp_bits_entry;
    end
    if (metaReset) begin
      _T_1038 <= 8'h0;
    end else if (io_bht_update_valid) begin
      if (io_bht_update_bits_branch) begin
        if (io_bht_update_bits_mispredict) begin
          _T_1038 <= _T_1121;
        end else if (io_bht_advance_valid) begin
          _T_1038 <= _T_1109;
        end
      end else if (io_bht_update_bits_mispredict) begin
        _T_1038 <= io_bht_update_bits_prediction_history;
      end else if (io_bht_advance_valid) begin
        _T_1038 <= _T_1109;
      end
    end else if (io_bht_advance_valid) begin
      _T_1038 <= _T_1109;
    end
    if (metaReset) begin
      _T_1125 <= 3'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1190) begin
        if (_T_1191) begin
          _T_1125 <= _T_1193;
        end
      end else if (_T_1199) begin
        if (~_T_1185) begin
          _T_1125 <= _T_1203;
        end
      end
    end
    if (metaReset) begin
      _T_1126 <= 3'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1190) begin
        if (_T_1194) begin
          _T_1126 <= _T_1197;
        end else begin
          _T_1126 <= 3'h0;
        end
      end else if (_T_1199) begin
        if (~_T_1185) begin
          if (_T_1204) begin
            _T_1126 <= _T_1207;
          end else begin
            _T_1126 <= 3'h5;
          end
        end
      end
    end
    if (metaReset) begin
      _T_1127_0 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1190) begin
        if (3'h0 == _T_1198) begin
          _T_1127_0 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      _T_1127_1 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1190) begin
        if (3'h1 == _T_1198) begin
          _T_1127_1 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      _T_1127_2 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1190) begin
        if (3'h2 == _T_1198) begin
          _T_1127_2 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      _T_1127_3 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1190) begin
        if (3'h3 == _T_1198) begin
          _T_1127_3 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      _T_1127_4 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1190) begin
        if (3'h4 == _T_1198) begin
          _T_1127_4 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      _T_1127_5 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1190) begin
        if (3'h5 == _T_1198) begin
          _T_1127_5 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    BTB_state <= BTB_xor0;
    if (!(BTB_cov_read_data)) begin
      BTB_covSum <= BTB_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(BTB_cov_write_en & BTB_cov_write_mask) begin
      BTB_cov[BTB_cov_write_addr] <= BTB_cov_write_data; // @[Coverage map for BTB]
    end
  end
endmodule
module TLMonitor_37(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [3:0]  io_in_a_bits_size,
  input  [1:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [7:0]  io_in_a_bits_mask,
  input         io_in_a_bits_corrupt,
  input         io_in_b_ready,
  input         io_in_b_valid,
  input  [2:0]  io_in_b_bits_opcode,
  input  [1:0]  io_in_b_bits_param,
  input  [3:0]  io_in_b_bits_size,
  input  [1:0]  io_in_b_bits_source,
  input  [31:0] io_in_b_bits_address,
  input  [7:0]  io_in_b_bits_mask,
  input         io_in_b_bits_corrupt,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [3:0]  io_in_c_bits_size,
  input  [1:0]  io_in_c_bits_source,
  input  [31:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [3:0]  io_in_d_bits_size,
  input  [1:0]  io_in_d_bits_source,
  input  [1:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_ready,
  input         io_in_e_valid,
  input  [1:0]  io_in_e_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire  _T_4; // @[Parameters.scala 47:9]
  wire  _T_5; // @[Parameters.scala 47:9]
  wire  _T_6; // @[Parameters.scala 47:9]
  wire  _T_8; // @[Parameters.scala 1016:46]
  wire  _T_9; // @[Parameters.scala 1016:46]
  wire [26:0] _T_11; // @[package.scala 212:77]
  wire [31:0] _GEN_71; // @[Edges.scala 22:16]
  wire [31:0] _T_14; // @[Edges.scala 22:16]
  wire  _T_15; // @[Edges.scala 22:24]
  wire [3:0] _T_18; // @[OneHot.scala 65:12]
  wire [2:0] _T_20; // @[Misc.scala 201:81]
  wire  _T_21; // @[Misc.scala 205:21]
  wire  _T_26; // @[Misc.scala 214:38]
  wire  _T_27; // @[Misc.scala 214:29]
  wire  _T_29; // @[Misc.scala 214:38]
  wire  _T_30; // @[Misc.scala 214:29]
  wire  _T_34; // @[Misc.scala 213:27]
  wire  _T_35; // @[Misc.scala 214:38]
  wire  _T_36; // @[Misc.scala 214:29]
  wire  _T_37; // @[Misc.scala 213:27]
  wire  _T_38; // @[Misc.scala 214:38]
  wire  _T_39; // @[Misc.scala 214:29]
  wire  _T_40; // @[Misc.scala 213:27]
  wire  _T_41; // @[Misc.scala 214:38]
  wire  _T_42; // @[Misc.scala 214:29]
  wire  _T_43; // @[Misc.scala 213:27]
  wire  _T_44; // @[Misc.scala 214:38]
  wire  _T_45; // @[Misc.scala 214:29]
  wire  _T_49; // @[Misc.scala 213:27]
  wire  _T_50; // @[Misc.scala 214:38]
  wire  _T_51; // @[Misc.scala 214:29]
  wire  _T_52; // @[Misc.scala 213:27]
  wire  _T_53; // @[Misc.scala 214:38]
  wire  _T_54; // @[Misc.scala 214:29]
  wire  _T_55; // @[Misc.scala 213:27]
  wire  _T_56; // @[Misc.scala 214:38]
  wire  _T_57; // @[Misc.scala 214:29]
  wire  _T_58; // @[Misc.scala 213:27]
  wire  _T_59; // @[Misc.scala 214:38]
  wire  _T_60; // @[Misc.scala 214:29]
  wire  _T_61; // @[Misc.scala 213:27]
  wire  _T_62; // @[Misc.scala 214:38]
  wire  _T_63; // @[Misc.scala 214:29]
  wire  _T_64; // @[Misc.scala 213:27]
  wire  _T_65; // @[Misc.scala 214:38]
  wire  _T_66; // @[Misc.scala 214:29]
  wire  _T_67; // @[Misc.scala 213:27]
  wire  _T_68; // @[Misc.scala 214:38]
  wire  _T_69; // @[Misc.scala 214:29]
  wire  _T_70; // @[Misc.scala 213:27]
  wire  _T_71; // @[Misc.scala 214:38]
  wire  _T_72; // @[Misc.scala 214:29]
  wire [7:0] _T_79; // @[Cat.scala 29:58]
  wire [32:0] _T_83; // @[Parameters.scala 137:49]
  wire  _T_109; // @[Monitor.scala 82:25]
  wire  _T_111; // @[Parameters.scala 93:42]
  wire  _T_118; // @[Parameters.scala 1066:30]
  wire  _T_128; // @[Parameters.scala 93:42]
  wire [31:0] _T_131; // @[Parameters.scala 137:31]
  wire [32:0] _T_132; // @[Parameters.scala 137:49]
  wire [32:0] _T_134; // @[Parameters.scala 137:52]
  wire  _T_135; // @[Parameters.scala 137:67]
  wire  _T_136; // @[Parameters.scala 601:56]
  wire  _T_139; // @[Parameters.scala 1240:195]
  wire  _T_141; // @[Monitor.scala 44:11]
  wire  _T_147; // @[Parameters.scala 92:48]
  wire  _T_148; // @[Mux.scala 27:72]
  wire  _T_165; // @[Parameters.scala 1255:195]
  wire  _T_167; // @[Monitor.scala 44:11]
  wire  _T_170; // @[Monitor.scala 44:11]
  wire  _T_174; // @[Monitor.scala 44:11]
  wire  _T_177; // @[Monitor.scala 44:11]
  wire  _T_179; // @[Bundles.scala 110:27]
  wire  _T_181; // @[Monitor.scala 44:11]
  wire  _T_184; // @[Monitor.scala 89:31]
  wire  _T_186; // @[Monitor.scala 44:11]
  wire  _T_190; // @[Monitor.scala 44:11]
  wire  _T_192; // @[Monitor.scala 93:25]
  wire  _T_266; // @[Monitor.scala 100:31]
  wire  _T_268; // @[Monitor.scala 44:11]
  wire  _T_279; // @[Monitor.scala 105:25]
  wire [31:0] _T_294; // @[Parameters.scala 137:31]
  wire [32:0] _T_295; // @[Parameters.scala 137:49]
  wire [32:0] _T_297; // @[Parameters.scala 137:52]
  wire  _T_298; // @[Parameters.scala 137:67]
  wire  _T_299; // @[Parameters.scala 601:56]
  wire [32:0] _T_307; // @[Parameters.scala 137:52]
  wire  _T_308; // @[Parameters.scala 137:67]
  wire [31:0] _T_309; // @[Parameters.scala 137:31]
  wire [32:0] _T_310; // @[Parameters.scala 137:49]
  wire [32:0] _T_312; // @[Parameters.scala 137:52]
  wire  _T_313; // @[Parameters.scala 137:67]
  wire [31:0] _T_314; // @[Parameters.scala 137:31]
  wire [32:0] _T_315; // @[Parameters.scala 137:49]
  wire [32:0] _T_317; // @[Parameters.scala 137:52]
  wire  _T_318; // @[Parameters.scala 137:67]
  wire [31:0] _T_319; // @[Parameters.scala 137:31]
  wire [32:0] _T_320; // @[Parameters.scala 137:49]
  wire [32:0] _T_322; // @[Parameters.scala 137:52]
  wire  _T_323; // @[Parameters.scala 137:67]
  wire [31:0] _T_324; // @[Parameters.scala 137:31]
  wire [32:0] _T_325; // @[Parameters.scala 137:49]
  wire [32:0] _T_327; // @[Parameters.scala 137:52]
  wire  _T_328; // @[Parameters.scala 137:67]
  wire [32:0] _T_332; // @[Parameters.scala 137:52]
  wire  _T_333; // @[Parameters.scala 137:67]
  wire  _T_334; // @[Parameters.scala 602:42]
  wire  _T_335; // @[Parameters.scala 602:42]
  wire  _T_336; // @[Parameters.scala 602:42]
  wire  _T_337; // @[Parameters.scala 602:42]
  wire  _T_338; // @[Parameters.scala 602:42]
  wire  _T_339; // @[Parameters.scala 601:56]
  wire  _T_341; // @[Parameters.scala 603:30]
  wire  _T_342; // @[Parameters.scala 1243:195]
  wire  _T_344; // @[Monitor.scala 44:11]
  wire  _T_352; // @[Monitor.scala 109:31]
  wire  _T_354; // @[Monitor.scala 44:11]
  wire  _T_356; // @[Monitor.scala 110:30]
  wire  _T_358; // @[Monitor.scala 44:11]
  wire  _T_364; // @[Monitor.scala 114:25]
  wire  _T_409; // @[Parameters.scala 602:42]
  wire  _T_410; // @[Parameters.scala 602:42]
  wire  _T_411; // @[Parameters.scala 602:42]
  wire  _T_412; // @[Parameters.scala 601:56]
  wire  _T_421; // @[Parameters.scala 93:42]
  wire  _T_429; // @[Parameters.scala 601:56]
  wire  _T_431; // @[Parameters.scala 603:30]
  wire  _T_433; // @[Parameters.scala 603:30]
  wire  _T_434; // @[Parameters.scala 1244:195]
  wire  _T_436; // @[Monitor.scala 44:11]
  wire  _T_452; // @[Monitor.scala 122:25]
  wire [7:0] _T_537; // @[Monitor.scala 127:31]
  wire  _T_538; // @[Monitor.scala 127:40]
  wire  _T_540; // @[Monitor.scala 44:11]
  wire  _T_542; // @[Monitor.scala 130:25]
  wire  _T_554; // @[Parameters.scala 93:42]
  wire [32:0] _T_560; // @[Parameters.scala 137:52]
  wire  _T_561; // @[Parameters.scala 137:67]
  wire  _T_567; // @[Parameters.scala 602:42]
  wire  _T_568; // @[Parameters.scala 601:56]
  wire  _T_590; // @[Parameters.scala 1241:195]
  wire  _T_592; // @[Monitor.scala 44:11]
  wire  _T_600; // @[Bundles.scala 140:33]
  wire  _T_602; // @[Monitor.scala 44:11]
  wire  _T_608; // @[Monitor.scala 138:25]
  wire  _T_666; // @[Bundles.scala 147:30]
  wire  _T_668; // @[Monitor.scala 44:11]
  wire  _T_674; // @[Monitor.scala 146:25]
  wire  _T_734; // @[Parameters.scala 1246:195]
  wire  _T_736; // @[Monitor.scala 44:11]
  wire  _T_744; // @[Bundles.scala 160:28]
  wire  _T_746; // @[Monitor.scala 44:11]
  wire  _T_756; // @[Bundles.scala 44:24]
  wire  _T_758; // @[Monitor.scala 51:11]
  wire  _T_760; // @[Parameters.scala 47:9]
  wire  _T_761; // @[Parameters.scala 47:9]
  wire  _T_762; // @[Parameters.scala 47:9]
  wire  _T_764; // @[Parameters.scala 1016:46]
  wire  _T_765; // @[Parameters.scala 1016:46]
  wire  _T_767; // @[Monitor.scala 310:25]
  wire  _T_769; // @[Monitor.scala 51:11]
  wire  _T_771; // @[Monitor.scala 312:27]
  wire  _T_773; // @[Monitor.scala 51:11]
  wire  _T_775; // @[Monitor.scala 313:28]
  wire  _T_777; // @[Monitor.scala 51:11]
  wire  _T_781; // @[Monitor.scala 51:11]
  wire  _T_785; // @[Monitor.scala 51:11]
  wire  _T_787; // @[Monitor.scala 318:25]
  wire  _T_798; // @[Bundles.scala 104:26]
  wire  _T_800; // @[Monitor.scala 51:11]
  wire  _T_802; // @[Monitor.scala 323:28]
  wire  _T_804; // @[Monitor.scala 51:11]
  wire  _T_815; // @[Monitor.scala 328:25]
  wire  _T_835; // @[Monitor.scala 334:30]
  wire  _T_837; // @[Monitor.scala 51:11]
  wire  _T_844; // @[Monitor.scala 338:25]
  wire  _T_861; // @[Monitor.scala 346:25]
  wire  _T_879; // @[Monitor.scala 354:25]
  wire  _T_896; // @[Bundles.scala 42:24]
  wire  _T_898; // @[Monitor.scala 44:11]
  wire  _T_900; // @[Parameters.scala 47:9]
  wire [32:0] _T_903; // @[Parameters.scala 137:49]
  wire  _T_908; // @[Parameters.scala 47:9]
  wire  _T_916; // @[Parameters.scala 47:9]
  wire [31:0] _T_929; // @[Parameters.scala 137:31]
  wire [32:0] _T_930; // @[Parameters.scala 137:49]
  wire [32:0] _T_932; // @[Parameters.scala 137:52]
  wire  _T_933; // @[Parameters.scala 137:67]
  wire [31:0] _T_934; // @[Parameters.scala 137:31]
  wire [32:0] _T_935; // @[Parameters.scala 137:49]
  wire [32:0] _T_937; // @[Parameters.scala 137:52]
  wire  _T_938; // @[Parameters.scala 137:67]
  wire [31:0] _T_939; // @[Parameters.scala 137:31]
  wire [32:0] _T_940; // @[Parameters.scala 137:49]
  wire [32:0] _T_942; // @[Parameters.scala 137:52]
  wire  _T_943; // @[Parameters.scala 137:67]
  wire [32:0] _T_947; // @[Parameters.scala 137:52]
  wire  _T_948; // @[Parameters.scala 137:67]
  wire [31:0] _T_949; // @[Parameters.scala 137:31]
  wire [32:0] _T_950; // @[Parameters.scala 137:49]
  wire [32:0] _T_952; // @[Parameters.scala 137:52]
  wire  _T_953; // @[Parameters.scala 137:67]
  wire [31:0] _T_954; // @[Parameters.scala 137:31]
  wire [32:0] _T_955; // @[Parameters.scala 137:49]
  wire [32:0] _T_957; // @[Parameters.scala 137:52]
  wire  _T_958; // @[Parameters.scala 137:67]
  wire [31:0] _T_959; // @[Parameters.scala 137:31]
  wire [32:0] _T_960; // @[Parameters.scala 137:49]
  wire [32:0] _T_962; // @[Parameters.scala 137:52]
  wire  _T_963; // @[Parameters.scala 137:67]
  wire  _T_965; // @[Parameters.scala 556:64]
  wire  _T_966; // @[Parameters.scala 556:64]
  wire  _T_967; // @[Parameters.scala 556:64]
  wire  _T_968; // @[Parameters.scala 556:64]
  wire  _T_969; // @[Parameters.scala 556:64]
  wire  _T_970; // @[Parameters.scala 556:64]
  wire [26:0] _T_972; // @[package.scala 212:77]
  wire [31:0] _GEN_72; // @[Edges.scala 22:16]
  wire [31:0] _T_975; // @[Edges.scala 22:16]
  wire  _T_976; // @[Edges.scala 22:24]
  wire [3:0] _T_979; // @[OneHot.scala 65:12]
  wire [2:0] _T_981; // @[Misc.scala 201:81]
  wire  _T_982; // @[Misc.scala 205:21]
  wire  _T_987; // @[Misc.scala 214:38]
  wire  _T_988; // @[Misc.scala 214:29]
  wire  _T_990; // @[Misc.scala 214:38]
  wire  _T_991; // @[Misc.scala 214:29]
  wire  _T_995; // @[Misc.scala 213:27]
  wire  _T_996; // @[Misc.scala 214:38]
  wire  _T_997; // @[Misc.scala 214:29]
  wire  _T_998; // @[Misc.scala 213:27]
  wire  _T_999; // @[Misc.scala 214:38]
  wire  _T_1000; // @[Misc.scala 214:29]
  wire  _T_1001; // @[Misc.scala 213:27]
  wire  _T_1002; // @[Misc.scala 214:38]
  wire  _T_1003; // @[Misc.scala 214:29]
  wire  _T_1004; // @[Misc.scala 213:27]
  wire  _T_1005; // @[Misc.scala 214:38]
  wire  _T_1006; // @[Misc.scala 214:29]
  wire  _T_1010; // @[Misc.scala 213:27]
  wire  _T_1011; // @[Misc.scala 214:38]
  wire  _T_1012; // @[Misc.scala 214:29]
  wire  _T_1013; // @[Misc.scala 213:27]
  wire  _T_1014; // @[Misc.scala 214:38]
  wire  _T_1015; // @[Misc.scala 214:29]
  wire  _T_1016; // @[Misc.scala 213:27]
  wire  _T_1017; // @[Misc.scala 214:38]
  wire  _T_1018; // @[Misc.scala 214:29]
  wire  _T_1019; // @[Misc.scala 213:27]
  wire  _T_1020; // @[Misc.scala 214:38]
  wire  _T_1021; // @[Misc.scala 214:29]
  wire  _T_1022; // @[Misc.scala 213:27]
  wire  _T_1023; // @[Misc.scala 214:38]
  wire  _T_1024; // @[Misc.scala 214:29]
  wire  _T_1025; // @[Misc.scala 213:27]
  wire  _T_1026; // @[Misc.scala 214:38]
  wire  _T_1027; // @[Misc.scala 214:29]
  wire  _T_1028; // @[Misc.scala 213:27]
  wire  _T_1029; // @[Misc.scala 214:38]
  wire  _T_1030; // @[Misc.scala 214:29]
  wire  _T_1031; // @[Misc.scala 213:27]
  wire  _T_1032; // @[Misc.scala 214:38]
  wire  _T_1033; // @[Misc.scala 214:29]
  wire [7:0] _T_1040; // @[Cat.scala 29:58]
  wire [1:0] _T_1047; // @[Mux.scala 27:72]
  wire [1:0] _GEN_73; // @[Mux.scala 27:72]
  wire [1:0] _T_1049; // @[Mux.scala 27:72]
  wire  _T_1051; // @[Monitor.scala 165:113]
  wire  _T_1052; // @[Monitor.scala 167:25]
  wire  _T_1057; // @[Parameters.scala 92:48]
  wire  _T_1058; // @[Mux.scala 27:72]
  wire  _T_1065; // @[Parameters.scala 93:42]
  wire  _T_1075; // @[Parameters.scala 1255:195]
  wire  _T_1077; // @[Monitor.scala 44:11]
  wire  _T_1080; // @[Monitor.scala 44:11]
  wire  _T_1083; // @[Monitor.scala 44:11]
  wire  _T_1086; // @[Monitor.scala 44:11]
  wire  _T_1088; // @[Bundles.scala 104:26]
  wire  _T_1090; // @[Monitor.scala 44:11]
  wire  _T_1092; // @[Monitor.scala 173:30]
  wire  _T_1094; // @[Monitor.scala 44:11]
  wire  _T_1098; // @[Monitor.scala 44:11]
  wire  _T_1100; // @[Monitor.scala 177:25]
  wire  _T_1125; // @[Monitor.scala 182:31]
  wire  _T_1127; // @[Monitor.scala 44:11]
  wire  _T_1137; // @[Monitor.scala 187:25]
  wire  _T_1170; // @[Monitor.scala 196:25]
  wire [7:0] _T_1200; // @[Monitor.scala 202:31]
  wire  _T_1201; // @[Monitor.scala 202:40]
  wire  _T_1203; // @[Monitor.scala 44:11]
  wire  _T_1205; // @[Monitor.scala 205:25]
  wire  _T_1238; // @[Monitor.scala 214:25]
  wire  _T_1271; // @[Monitor.scala 223:25]
  wire  _T_1308; // @[Parameters.scala 47:9]
  wire  _T_1309; // @[Parameters.scala 47:9]
  wire  _T_1310; // @[Parameters.scala 47:9]
  wire  _T_1312; // @[Parameters.scala 1016:46]
  wire  _T_1313; // @[Parameters.scala 1016:46]
  wire [26:0] _T_1315; // @[package.scala 212:77]
  wire [31:0] _GEN_74; // @[Edges.scala 22:16]
  wire [31:0] _T_1318; // @[Edges.scala 22:16]
  wire  _T_1319; // @[Edges.scala 22:24]
  wire [31:0] _T_1320; // @[Parameters.scala 137:31]
  wire [32:0] _T_1321; // @[Parameters.scala 137:49]
  wire [32:0] _T_1323; // @[Parameters.scala 137:52]
  wire  _T_1324; // @[Parameters.scala 137:67]
  wire [31:0] _T_1325; // @[Parameters.scala 137:31]
  wire [32:0] _T_1326; // @[Parameters.scala 137:49]
  wire [32:0] _T_1328; // @[Parameters.scala 137:52]
  wire  _T_1329; // @[Parameters.scala 137:67]
  wire [31:0] _T_1330; // @[Parameters.scala 137:31]
  wire [32:0] _T_1331; // @[Parameters.scala 137:49]
  wire [32:0] _T_1333; // @[Parameters.scala 137:52]
  wire  _T_1334; // @[Parameters.scala 137:67]
  wire [32:0] _T_1336; // @[Parameters.scala 137:49]
  wire [32:0] _T_1338; // @[Parameters.scala 137:52]
  wire  _T_1339; // @[Parameters.scala 137:67]
  wire [31:0] _T_1340; // @[Parameters.scala 137:31]
  wire [32:0] _T_1341; // @[Parameters.scala 137:49]
  wire [32:0] _T_1343; // @[Parameters.scala 137:52]
  wire  _T_1344; // @[Parameters.scala 137:67]
  wire [31:0] _T_1345; // @[Parameters.scala 137:31]
  wire [32:0] _T_1346; // @[Parameters.scala 137:49]
  wire [32:0] _T_1348; // @[Parameters.scala 137:52]
  wire  _T_1349; // @[Parameters.scala 137:67]
  wire [31:0] _T_1350; // @[Parameters.scala 137:31]
  wire [32:0] _T_1351; // @[Parameters.scala 137:49]
  wire [32:0] _T_1353; // @[Parameters.scala 137:52]
  wire  _T_1354; // @[Parameters.scala 137:67]
  wire  _T_1356; // @[Parameters.scala 556:64]
  wire  _T_1357; // @[Parameters.scala 556:64]
  wire  _T_1358; // @[Parameters.scala 556:64]
  wire  _T_1359; // @[Parameters.scala 556:64]
  wire  _T_1360; // @[Parameters.scala 556:64]
  wire  _T_1361; // @[Parameters.scala 556:64]
  wire  _T_1391; // @[Monitor.scala 242:25]
  wire  _T_1393; // @[Monitor.scala 44:11]
  wire  _T_1396; // @[Monitor.scala 44:11]
  wire  _T_1398; // @[Monitor.scala 245:30]
  wire  _T_1400; // @[Monitor.scala 44:11]
  wire  _T_1403; // @[Monitor.scala 44:11]
  wire  _T_1405; // @[Bundles.scala 122:29]
  wire  _T_1407; // @[Monitor.scala 44:11]
  wire  _T_1413; // @[Monitor.scala 251:25]
  wire  _T_1431; // @[Monitor.scala 259:25]
  wire  _T_1433; // @[Parameters.scala 93:42]
  wire  _T_1440; // @[Parameters.scala 1066:30]
  wire  _T_1450; // @[Parameters.scala 93:42]
  wire [32:0] _T_1456; // @[Parameters.scala 137:52]
  wire  _T_1457; // @[Parameters.scala 137:67]
  wire  _T_1458; // @[Parameters.scala 601:56]
  wire  _T_1461; // @[Parameters.scala 1240:195]
  wire  _T_1463; // @[Monitor.scala 44:11]
  wire  _T_1469; // @[Parameters.scala 92:48]
  wire  _T_1470; // @[Mux.scala 27:72]
  wire  _T_1487; // @[Parameters.scala 1255:195]
  wire  _T_1489; // @[Monitor.scala 44:11]
  wire  _T_1501; // @[Bundles.scala 116:29]
  wire  _T_1503; // @[Monitor.scala 44:11]
  wire  _T_1509; // @[Monitor.scala 269:25]
  wire  _T_1583; // @[Monitor.scala 278:25]
  wire  _T_1593; // @[Monitor.scala 282:31]
  wire  _T_1595; // @[Monitor.scala 44:11]
  wire  _T_1601; // @[Monitor.scala 286:25]
  wire  _T_1615; // @[Monitor.scala 293:25]
  wire  _T_1637; // @[Decoupled.scala 40:37]
  wire [8:0] _T_1642; // @[Edges.scala 221:59]
  reg [8:0] _T_1646; // @[Edges.scala 230:27]
  reg [31:0] _RAND_0;
  wire [8:0] _T_1648; // @[Edges.scala 231:28]
  wire  _T_1649; // @[Edges.scala 232:25]
  reg [2:0] _T_1657; // @[Monitor.scala 384:22]
  reg [31:0] _RAND_1;
  reg [2:0] _T_1658; // @[Monitor.scala 385:22]
  reg [31:0] _RAND_2;
  reg [3:0] _T_1659; // @[Monitor.scala 386:22]
  reg [31:0] _RAND_3;
  reg [1:0] _T_1660; // @[Monitor.scala 387:22]
  reg [31:0] _RAND_4;
  reg [31:0] _T_1661; // @[Monitor.scala 388:22]
  reg [31:0] _RAND_5;
  wire  _T_1663; // @[Monitor.scala 389:19]
  wire  _T_1664; // @[Monitor.scala 390:32]
  wire  _T_1666; // @[Monitor.scala 44:11]
  wire  _T_1668; // @[Monitor.scala 391:32]
  wire  _T_1670; // @[Monitor.scala 44:11]
  wire  _T_1672; // @[Monitor.scala 392:32]
  wire  _T_1674; // @[Monitor.scala 44:11]
  wire  _T_1676; // @[Monitor.scala 393:32]
  wire  _T_1678; // @[Monitor.scala 44:11]
  wire  _T_1680; // @[Monitor.scala 394:32]
  wire  _T_1682; // @[Monitor.scala 44:11]
  wire  _T_1685; // @[Monitor.scala 396:20]
  wire  _T_1686; // @[Decoupled.scala 40:37]
  wire [26:0] _T_1688; // @[package.scala 212:77]
  wire [8:0] _T_1691; // @[Edges.scala 221:59]
  reg [8:0] _T_1694; // @[Edges.scala 230:27]
  reg [31:0] _RAND_6;
  wire [8:0] _T_1696; // @[Edges.scala 231:28]
  wire  _T_1697; // @[Edges.scala 232:25]
  reg [2:0] _T_1705; // @[Monitor.scala 535:22]
  reg [31:0] _RAND_7;
  reg [1:0] _T_1706; // @[Monitor.scala 536:22]
  reg [31:0] _RAND_8;
  reg [3:0] _T_1707; // @[Monitor.scala 537:22]
  reg [31:0] _RAND_9;
  reg [1:0] _T_1708; // @[Monitor.scala 538:22]
  reg [31:0] _RAND_10;
  reg [1:0] _T_1709; // @[Monitor.scala 539:22]
  reg [31:0] _RAND_11;
  reg  _T_1710; // @[Monitor.scala 540:22]
  reg [31:0] _RAND_12;
  wire  _T_1712; // @[Monitor.scala 541:19]
  wire  _T_1713; // @[Monitor.scala 542:29]
  wire  _T_1715; // @[Monitor.scala 51:11]
  wire  _T_1717; // @[Monitor.scala 543:29]
  wire  _T_1719; // @[Monitor.scala 51:11]
  wire  _T_1721; // @[Monitor.scala 544:29]
  wire  _T_1723; // @[Monitor.scala 51:11]
  wire  _T_1725; // @[Monitor.scala 545:29]
  wire  _T_1727; // @[Monitor.scala 51:11]
  wire  _T_1729; // @[Monitor.scala 546:29]
  wire  _T_1731; // @[Monitor.scala 51:11]
  wire  _T_1733; // @[Monitor.scala 547:29]
  wire  _T_1735; // @[Monitor.scala 51:11]
  wire  _T_1738; // @[Monitor.scala 549:20]
  wire  _T_1739; // @[Decoupled.scala 40:37]
  reg [8:0] _T_1748; // @[Edges.scala 230:27]
  reg [31:0] _RAND_13;
  wire [8:0] _T_1750; // @[Edges.scala 231:28]
  wire  _T_1751; // @[Edges.scala 232:25]
  reg [2:0] _T_1759; // @[Monitor.scala 407:22]
  reg [31:0] _RAND_14;
  reg [1:0] _T_1760; // @[Monitor.scala 408:22]
  reg [31:0] _RAND_15;
  reg [3:0] _T_1761; // @[Monitor.scala 409:22]
  reg [31:0] _RAND_16;
  reg [1:0] _T_1762; // @[Monitor.scala 410:22]
  reg [31:0] _RAND_17;
  reg [31:0] _T_1763; // @[Monitor.scala 411:22]
  reg [31:0] _RAND_18;
  wire  _T_1765; // @[Monitor.scala 412:19]
  wire  _T_1766; // @[Monitor.scala 413:32]
  wire  _T_1768; // @[Monitor.scala 44:11]
  wire  _T_1770; // @[Monitor.scala 414:32]
  wire  _T_1772; // @[Monitor.scala 44:11]
  wire  _T_1774; // @[Monitor.scala 415:32]
  wire  _T_1776; // @[Monitor.scala 44:11]
  wire  _T_1778; // @[Monitor.scala 416:32]
  wire  _T_1780; // @[Monitor.scala 44:11]
  wire  _T_1782; // @[Monitor.scala 417:32]
  wire  _T_1784; // @[Monitor.scala 44:11]
  wire  _T_1787; // @[Monitor.scala 419:20]
  wire  _T_1788; // @[Decoupled.scala 40:37]
  wire [8:0] _T_1793; // @[Edges.scala 221:59]
  reg [8:0] _T_1796; // @[Edges.scala 230:27]
  reg [31:0] _RAND_19;
  wire [8:0] _T_1798; // @[Edges.scala 231:28]
  wire  _T_1799; // @[Edges.scala 232:25]
  reg [2:0] _T_1807; // @[Monitor.scala 512:22]
  reg [31:0] _RAND_20;
  reg [2:0] _T_1808; // @[Monitor.scala 513:22]
  reg [31:0] _RAND_21;
  reg [3:0] _T_1809; // @[Monitor.scala 514:22]
  reg [31:0] _RAND_22;
  reg [1:0] _T_1810; // @[Monitor.scala 515:22]
  reg [31:0] _RAND_23;
  reg [31:0] _T_1811; // @[Monitor.scala 516:22]
  reg [31:0] _RAND_24;
  wire  _T_1813; // @[Monitor.scala 517:19]
  wire  _T_1814; // @[Monitor.scala 518:32]
  wire  _T_1816; // @[Monitor.scala 44:11]
  wire  _T_1818; // @[Monitor.scala 519:32]
  wire  _T_1820; // @[Monitor.scala 44:11]
  wire  _T_1822; // @[Monitor.scala 520:32]
  wire  _T_1824; // @[Monitor.scala 44:11]
  wire  _T_1826; // @[Monitor.scala 521:32]
  wire  _T_1828; // @[Monitor.scala 44:11]
  wire  _T_1830; // @[Monitor.scala 522:32]
  wire  _T_1832; // @[Monitor.scala 44:11]
  wire  _T_1835; // @[Monitor.scala 524:20]
  reg [2:0] inflight; // @[Monitor.scala 611:27]
  reg [31:0] _RAND_25;
  reg [11:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [31:0] _RAND_26;
  reg [23:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [31:0] _RAND_27;
  reg [8:0] _T_1845; // @[Edges.scala 230:27]
  reg [31:0] _RAND_28;
  wire [8:0] _T_1847; // @[Edges.scala 231:28]
  wire  a_first; // @[Edges.scala 232:25]
  reg [8:0] _T_1863; // @[Edges.scala 230:27]
  reg [31:0] _RAND_29;
  wire [8:0] _T_1865; // @[Edges.scala 231:28]
  wire  d_first; // @[Edges.scala 232:25]
  wire [3:0] _GEN_75; // @[Monitor.scala 632:69]
  wire [4:0] _T_1873; // @[Monitor.scala 632:69]
  wire [11:0] _T_1874; // @[Monitor.scala 632:44]
  wire [15:0] _T_1878; // @[Monitor.scala 609:57]
  wire [15:0] _GEN_76; // @[Monitor.scala 632:97]
  wire [15:0] _T_1879; // @[Monitor.scala 632:97]
  wire [15:0] _T_1880; // @[Monitor.scala 632:152]
  wire [4:0] _T_1881; // @[Monitor.scala 636:65]
  wire [23:0] _T_1882; // @[Monitor.scala 636:40]
  wire [15:0] _T_1886; // @[Monitor.scala 609:57]
  wire [23:0] _GEN_78; // @[Monitor.scala 636:91]
  wire [23:0] _T_1887; // @[Monitor.scala 636:91]
  wire [23:0] _T_1888; // @[Monitor.scala 636:144]
  wire  _T_1892; // @[Monitor.scala 646:27]
  wire [3:0] _T_1894; // @[OneHot.scala 58:35]
  wire [3:0] _T_1895; // @[Monitor.scala 648:53]
  wire [3:0] _T_1896; // @[Monitor.scala 648:61]
  wire [4:0] _T_1897; // @[Monitor.scala 649:49]
  wire [4:0] _T_1898; // @[Monitor.scala 649:57]
  wire [3:0] _GEN_80; // @[Monitor.scala 650:72]
  wire [4:0] _T_1899; // @[Monitor.scala 650:72]
  wire [3:0] a_opcodes_set_interm; // @[Monitor.scala 646:72]
  wire [34:0] _GEN_81; // @[Monitor.scala 650:47]
  wire [34:0] _T_1900; // @[Monitor.scala 650:47]
  wire [4:0] _T_1901; // @[Monitor.scala 651:68]
  wire [4:0] a_sizes_set_interm; // @[Monitor.scala 646:72]
  wire [35:0] _GEN_82; // @[Monitor.scala 651:43]
  wire [35:0] _T_1902; // @[Monitor.scala 651:43]
  wire [2:0] _T_1903; // @[Monitor.scala 652:26]
  wire  _T_1907; // @[Monitor.scala 44:11]
  wire [3:0] _GEN_27; // @[Monitor.scala 646:72]
  wire [34:0] _GEN_30; // @[Monitor.scala 646:72]
  wire [35:0] _GEN_31; // @[Monitor.scala 646:72]
  wire  _T_1911; // @[Monitor.scala 663:27]
  wire  _T_1914; // @[Monitor.scala 663:72]
  wire [3:0] _T_1915; // @[OneHot.scala 58:35]
  wire [46:0] _GEN_84; // @[Monitor.scala 665:76]
  wire [46:0] _T_1921; // @[Monitor.scala 665:76]
  wire [46:0] _GEN_85; // @[Monitor.scala 666:72]
  wire [46:0] _T_1927; // @[Monitor.scala 666:72]
  wire [3:0] _GEN_32; // @[Monitor.scala 663:91]
  wire [46:0] _GEN_33; // @[Monitor.scala 663:91]
  wire [46:0] _GEN_34; // @[Monitor.scala 663:91]
  wire  _T_1928; // @[Monitor.scala 668:26]
  wire  _T_1931; // @[Monitor.scala 668:71]
  wire [2:0] _T_1932; // @[Monitor.scala 669:25]
  wire  _T_1934; // @[Monitor.scala 669:93]
  wire  _T_1935; // @[Monitor.scala 669:68]
  wire  _T_1936; // @[Monitor.scala 669:142]
  wire  _T_1937; // @[Monitor.scala 669:119]
  wire  _T_1938; // @[Monitor.scala 669:166]
  wire  _T_1939; // @[Monitor.scala 669:49]
  wire  _T_1941; // @[Monitor.scala 51:11]
  wire [3:0] a_opcode_lookup; // @[Monitor.scala 632:21]
  wire [2:0] _GEN_37; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_38; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_39; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_40; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_41; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_42; // @[Monitor.scala 670:37]
  wire  _T_1944; // @[Monitor.scala 670:37]
  wire [2:0] _GEN_49; // @[Monitor.scala 670:96]
  wire [2:0] _GEN_50; // @[Monitor.scala 670:96]
  wire  _T_1946; // @[Monitor.scala 670:96]
  wire  _T_1947; // @[Monitor.scala 670:71]
  wire [2:0] _GEN_53; // @[Monitor.scala 671:60]
  wire [2:0] _GEN_54; // @[Monitor.scala 671:60]
  wire [2:0] _GEN_55; // @[Monitor.scala 671:60]
  wire [2:0] _GEN_56; // @[Monitor.scala 671:60]
  wire [2:0] _GEN_57; // @[Monitor.scala 671:60]
  wire [2:0] _GEN_58; // @[Monitor.scala 671:60]
  wire  _T_1948; // @[Monitor.scala 671:60]
  wire [2:0] _GEN_65; // @[Monitor.scala 671:124]
  wire [2:0] _GEN_66; // @[Monitor.scala 671:124]
  wire  _T_1949; // @[Monitor.scala 671:124]
  wire  _T_1950; // @[Monitor.scala 671:99]
  wire  _T_1951; // @[Monitor.scala 671:34]
  wire  _T_1952; // @[Monitor.scala 671:15]
  wire  _T_1954; // @[Monitor.scala 51:11]
  wire [7:0] a_size_lookup; // @[Monitor.scala 636:19]
  wire [7:0] _GEN_86; // @[Monitor.scala 673:34]
  wire  _T_1956; // @[Monitor.scala 673:34]
  wire  _T_1958; // @[Monitor.scala 673:72]
  wire  _T_1959; // @[Monitor.scala 673:53]
  wire  _T_1961; // @[Monitor.scala 51:11]
  wire  _T_1964; // @[Monitor.scala 675:36]
  wire  _T_1965; // @[Monitor.scala 675:47]
  wire  _T_1967; // @[Monitor.scala 675:65]
  wire  _T_1969; // @[Monitor.scala 675:116]
  wire  _T_1971; // @[Monitor.scala 676:32]
  wire  _T_1973; // @[Monitor.scala 51:11]
  wire [2:0] a_set; // @[Monitor.scala 647:13]
  wire [2:0] d_clr; // @[Monitor.scala 664:13]
  wire  _T_1975; // @[Monitor.scala 680:20]
  wire  _T_1976; // @[Monitor.scala 680:40]
  wire  _T_1978; // @[Monitor.scala 680:30]
  wire  _T_1980; // @[Monitor.scala 51:11]
  wire [2:0] _T_1982; // @[Monitor.scala 683:27]
  wire [2:0] _T_1984; // @[Monitor.scala 683:36]
  wire [11:0] a_opcodes_set; // @[Monitor.scala 650:21]
  wire [11:0] _T_1985; // @[Monitor.scala 684:43]
  wire [11:0] d_opcodes_clr; // @[Monitor.scala 665:21]
  wire [11:0] _T_1987; // @[Monitor.scala 684:60]
  wire [23:0] a_sizes_set; // @[Monitor.scala 651:19]
  wire [23:0] _T_1988; // @[Monitor.scala 685:39]
  wire [23:0] d_sizes_clr; // @[Monitor.scala 666:19]
  wire [23:0] _T_1990; // @[Monitor.scala 685:54]
  reg [3:0] _T_2006; // @[Monitor.scala 697:27]
  reg [31:0] _RAND_30;
  reg [8:0] _T_2015; // @[Edges.scala 230:27]
  reg [31:0] _RAND_31;
  wire [8:0] _T_2017; // @[Edges.scala 231:28]
  wire  _T_2018; // @[Edges.scala 232:25]
  wire  _T_2028; // @[Monitor.scala 703:27]
  wire  _T_2032; // @[Edges.scala 72:40]
  wire  _T_2033; // @[Monitor.scala 703:38]
  wire [3:0] _T_2034; // @[OneHot.scala 58:35]
  wire [3:0] _T_2035; // @[Monitor.scala 705:23]
  wire  _T_2039; // @[Monitor.scala 51:11]
  wire [3:0] _GEN_69; // @[Monitor.scala 703:72]
  wire  _T_2042; // @[Decoupled.scala 40:37]
  wire [3:0] _T_2045; // @[OneHot.scala 58:35]
  wire [3:0] _T_2046; // @[Monitor.scala 711:24]
  wire [3:0] _T_2047; // @[Monitor.scala 711:35]
  wire  _T_2050; // @[Monitor.scala 44:11]
  wire [3:0] _GEN_70; // @[Monitor.scala 709:73]
  wire [3:0] _T_2052; // @[Monitor.scala 716:27]
  wire [3:0] _T_2054; // @[Monitor.scala 716:36]
  wire  _GEN_87; // @[Monitor.scala 44:11]
  wire  _GEN_103; // @[Monitor.scala 44:11]
  wire  _GEN_121; // @[Monitor.scala 44:11]
  wire  _GEN_133; // @[Monitor.scala 44:11]
  wire  _GEN_143; // @[Monitor.scala 44:11]
  wire  _GEN_153; // @[Monitor.scala 44:11]
  wire  _GEN_163; // @[Monitor.scala 44:11]
  wire  _GEN_173; // @[Monitor.scala 44:11]
  wire  _GEN_185; // @[Monitor.scala 51:11]
  wire  _GEN_195; // @[Monitor.scala 51:11]
  wire  _GEN_205; // @[Monitor.scala 51:11]
  wire  _GEN_215; // @[Monitor.scala 51:11]
  wire  _GEN_221; // @[Monitor.scala 51:11]
  wire  _GEN_227; // @[Monitor.scala 51:11]
  wire  _GEN_233; // @[Monitor.scala 44:11]
  wire  _GEN_247; // @[Monitor.scala 44:11]
  wire  _GEN_261; // @[Monitor.scala 44:11]
  wire  _GEN_273; // @[Monitor.scala 44:11]
  wire  _GEN_285; // @[Monitor.scala 44:11]
  wire  _GEN_295; // @[Monitor.scala 44:11]
  wire  _GEN_305; // @[Monitor.scala 44:11]
  wire  _GEN_317; // @[Monitor.scala 44:11]
  wire  _GEN_327; // @[Monitor.scala 44:11]
  wire  _GEN_337; // @[Monitor.scala 44:11]
  wire  _GEN_349; // @[Monitor.scala 44:11]
  wire  _GEN_361; // @[Monitor.scala 44:11]
  wire  _GEN_369; // @[Monitor.scala 44:11]
  wire  _GEN_377; // @[Monitor.scala 44:11]
  wire [29:0] TLMonitor_37_covSum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  stopEn4;
  wire  stopEn5;
  wire  stopEn6;
  wire  stopEn7;
  wire  stopEn8;
  wire  stopEn9;
  wire  stopEn10;
  wire  stopEn11;
  wire  stopEn12;
  wire  stopEn13;
  wire  stopEn14;
  wire  stopEn15;
  wire  stopEn16;
  wire  stopEn17;
  wire  stopEn18;
  wire  stopEn19;
  wire  stopEn20;
  wire  stopEn21;
  wire  stopEn22;
  wire  stopEn23;
  wire  stopEn24;
  wire  stopEn25;
  wire  stopEn26;
  wire  stopEn27;
  wire  stopEn28;
  wire  stopEn29;
  wire  stopEn30;
  wire  stopEn31;
  wire  stopEn32;
  wire  stopEn33;
  wire  stopEn34;
  wire  stopEn35;
  wire  stopEn36;
  wire  stopEn37;
  wire  stopEn38;
  wire  stopEn39;
  wire  stopEn40;
  wire  stopEn41;
  wire  stopEn42;
  wire  stopEn43;
  wire  stopEn44;
  wire  stopEn45;
  wire  stopEn46;
  wire  stopEn47;
  wire  stopEn48;
  wire  stopEn49;
  wire  stopEn50;
  wire  stopEn51;
  wire  stopEn52;
  wire  stopEn53;
  wire  stopEn54;
  wire  stopEn55;
  wire  stopEn56;
  wire  stopEn57;
  wire  stopEn58;
  wire  stopEn59;
  wire  stopEn60;
  wire  stopEn61;
  wire  stopEn62;
  wire  stopEn63;
  wire  stopEn64;
  wire  stopEn65;
  wire  stopEn66;
  wire  stopEn67;
  wire  stopEn68;
  wire  stopEn69;
  wire  stopEn70;
  wire  stopEn71;
  wire  stopEn72;
  wire  stopEn73;
  wire  stopEn74;
  wire  stopEn75;
  wire  stopEn76;
  wire  stopEn77;
  wire  stopEn78;
  wire  stopEn79;
  wire  stopEn80;
  wire  stopEn81;
  wire  stopEn82;
  wire  stopEn83;
  wire  stopEn84;
  wire  stopEn85;
  wire  stopEn86;
  wire  stopEn87;
  wire  stopEn88;
  wire  stopEn89;
  wire  stopEn90;
  wire  stopEn91;
  wire  stopEn92;
  wire  stopEn93;
  wire  stopEn94;
  wire  stopEn95;
  wire  stopEn96;
  wire  stopEn97;
  wire  stopEn98;
  wire  stopEn99;
  wire  stopEn100;
  wire  stopEn101;
  wire  stopEn102;
  wire  stopEn103;
  wire  stopEn104;
  wire  stopEn105;
  wire  stopEn106;
  wire  stopEn107;
  wire  stopEn108;
  wire  stopEn109;
  wire  stopEn110;
  wire  stopEn111;
  wire  stopEn112;
  wire  stopEn113;
  wire  stopEn114;
  wire  stopEn115;
  wire  stopEn116;
  wire  stopEn117;
  wire  stopEn118;
  wire  stopEn119;
  wire  stopEn120;
  wire  stopEn121;
  wire  stopEn122;
  wire  stopEn123;
  wire  stopEn124;
  wire  stopEn125;
  wire  stopEn126;
  wire  stopEn127;
  wire  stopEn128;
  wire  stopEn129;
  wire  stopEn130;
  wire  stopEn131;
  wire  stopEn132;
  wire  stopEn133;
  wire  stopEn134;
  wire  stopEn135;
  wire  stopEn136;
  wire  stopEn137;
  wire  stopEn138;
  wire  stopEn139;
  wire  stopEn140;
  wire  stopEn141;
  wire  stopEn142;
  wire  stopEn143;
  wire  stopEn144;
  wire  stopEn145;
  wire  stopEn146;
  wire  stopEn147;
  wire  stopEn148;
  wire  stopEn149;
  wire  stopEn150;
  wire  stopEn151;
  wire  stopEn152;
  wire  stopEn153;
  wire  stopEn154;
  wire  stopEn155;
  wire  stopEn156;
  wire  stopEn157;
  wire  stopEn158;
  wire  stopEn159;
  wire  stopEn160;
  wire  stopEn161;
  wire  stopEn162;
  wire  stopEn163;
  wire  stopEn164;
  wire  stopEn165;
  wire  stopEn166;
  wire  stopEn167;
  wire  stopEn168;
  wire  stopEn169;
  wire  stopEn170;
  wire  stopEn171;
  wire  stopEn172;
  wire  stopEn173;
  wire  stopEn174;
  wire  stopEn175;
  wire  stopEn176;
  wire  stopEn177;
  wire  stopEn178;
  wire  stopEn179;
  wire  TLMonitor_37_or63;
  wire  TLMonitor_37_or130;
  wire  TLMonitor_37_or64;
  wire  TLMonitor_37_or31;
  wire  TLMonitor_37_or132;
  wire  TLMonitor_37_or65;
  wire  TLMonitor_37_or134;
  wire  TLMonitor_37_or66;
  wire  TLMonitor_37_or32;
  wire  TLMonitor_37_or15;
  wire  TLMonitor_37_or67;
  wire  TLMonitor_37_or138;
  wire  TLMonitor_37_or68;
  wire  TLMonitor_37_or33;
  wire  TLMonitor_37_or140;
  wire  TLMonitor_37_or69;
  wire  TLMonitor_37_or142;
  wire  TLMonitor_37_or70;
  wire  TLMonitor_37_or34;
  wire  TLMonitor_37_or16;
  wire  TLMonitor_37_or7;
  wire  TLMonitor_37_or71;
  wire  TLMonitor_37_or146;
  wire  TLMonitor_37_or72;
  wire  TLMonitor_37_or35;
  wire  TLMonitor_37_or148;
  wire  TLMonitor_37_or73;
  wire  TLMonitor_37_or150;
  wire  TLMonitor_37_or74;
  wire  TLMonitor_37_or36;
  wire  TLMonitor_37_or17;
  wire  TLMonitor_37_or152;
  wire  TLMonitor_37_or75;
  wire  TLMonitor_37_or154;
  wire  TLMonitor_37_or76;
  wire  TLMonitor_37_or37;
  wire  TLMonitor_37_or156;
  wire  TLMonitor_37_or77;
  wire  TLMonitor_37_or158;
  wire  TLMonitor_37_or78;
  wire  TLMonitor_37_or38;
  wire  TLMonitor_37_or18;
  wire  TLMonitor_37_or8;
  wire  TLMonitor_37_or3;
  wire  TLMonitor_37_or79;
  wire  TLMonitor_37_or162;
  wire  TLMonitor_37_or80;
  wire  TLMonitor_37_or39;
  wire  TLMonitor_37_or164;
  wire  TLMonitor_37_or81;
  wire  TLMonitor_37_or166;
  wire  TLMonitor_37_or82;
  wire  TLMonitor_37_or40;
  wire  TLMonitor_37_or19;
  wire  TLMonitor_37_or83;
  wire  TLMonitor_37_or170;
  wire  TLMonitor_37_or84;
  wire  TLMonitor_37_or41;
  wire  TLMonitor_37_or172;
  wire  TLMonitor_37_or85;
  wire  TLMonitor_37_or174;
  wire  TLMonitor_37_or86;
  wire  TLMonitor_37_or42;
  wire  TLMonitor_37_or20;
  wire  TLMonitor_37_or9;
  wire  TLMonitor_37_or87;
  wire  TLMonitor_37_or178;
  wire  TLMonitor_37_or88;
  wire  TLMonitor_37_or43;
  wire  TLMonitor_37_or180;
  wire  TLMonitor_37_or89;
  wire  TLMonitor_37_or182;
  wire  TLMonitor_37_or90;
  wire  TLMonitor_37_or44;
  wire  TLMonitor_37_or21;
  wire  TLMonitor_37_or184;
  wire  TLMonitor_37_or91;
  wire  TLMonitor_37_or186;
  wire  TLMonitor_37_or92;
  wire  TLMonitor_37_or45;
  wire  TLMonitor_37_or188;
  wire  TLMonitor_37_or93;
  wire  TLMonitor_37_or190;
  wire  TLMonitor_37_or94;
  wire  TLMonitor_37_or46;
  wire  TLMonitor_37_or22;
  wire  TLMonitor_37_or10;
  wire  TLMonitor_37_or4;
  wire  TLMonitor_37_or1;
  wire  TLMonitor_37_or95;
  wire  TLMonitor_37_or194;
  wire  TLMonitor_37_or96;
  wire  TLMonitor_37_or47;
  wire  TLMonitor_37_or196;
  wire  TLMonitor_37_or97;
  wire  TLMonitor_37_or198;
  wire  TLMonitor_37_or98;
  wire  TLMonitor_37_or48;
  wire  TLMonitor_37_or23;
  wire  TLMonitor_37_or99;
  wire  TLMonitor_37_or202;
  wire  TLMonitor_37_or100;
  wire  TLMonitor_37_or49;
  wire  TLMonitor_37_or204;
  wire  TLMonitor_37_or101;
  wire  TLMonitor_37_or206;
  wire  TLMonitor_37_or102;
  wire  TLMonitor_37_or50;
  wire  TLMonitor_37_or24;
  wire  TLMonitor_37_or11;
  wire  TLMonitor_37_or103;
  wire  TLMonitor_37_or210;
  wire  TLMonitor_37_or104;
  wire  TLMonitor_37_or51;
  wire  TLMonitor_37_or212;
  wire  TLMonitor_37_or105;
  wire  TLMonitor_37_or214;
  wire  TLMonitor_37_or106;
  wire  TLMonitor_37_or52;
  wire  TLMonitor_37_or25;
  wire  TLMonitor_37_or216;
  wire  TLMonitor_37_or107;
  wire  TLMonitor_37_or218;
  wire  TLMonitor_37_or108;
  wire  TLMonitor_37_or53;
  wire  TLMonitor_37_or220;
  wire  TLMonitor_37_or109;
  wire  TLMonitor_37_or222;
  wire  TLMonitor_37_or110;
  wire  TLMonitor_37_or54;
  wire  TLMonitor_37_or26;
  wire  TLMonitor_37_or12;
  wire  TLMonitor_37_or5;
  wire  TLMonitor_37_or111;
  wire  TLMonitor_37_or226;
  wire  TLMonitor_37_or112;
  wire  TLMonitor_37_or55;
  wire  TLMonitor_37_or228;
  wire  TLMonitor_37_or113;
  wire  TLMonitor_37_or230;
  wire  TLMonitor_37_or114;
  wire  TLMonitor_37_or56;
  wire  TLMonitor_37_or27;
  wire  TLMonitor_37_or115;
  wire  TLMonitor_37_or234;
  wire  TLMonitor_37_or116;
  wire  TLMonitor_37_or57;
  wire  TLMonitor_37_or236;
  wire  TLMonitor_37_or117;
  wire  TLMonitor_37_or238;
  wire  TLMonitor_37_or118;
  wire  TLMonitor_37_or58;
  wire  TLMonitor_37_or28;
  wire  TLMonitor_37_or13;
  wire  TLMonitor_37_or119;
  wire  TLMonitor_37_or242;
  wire  TLMonitor_37_or120;
  wire  TLMonitor_37_or59;
  wire  TLMonitor_37_or244;
  wire  TLMonitor_37_or121;
  wire  TLMonitor_37_or246;
  wire  TLMonitor_37_or122;
  wire  TLMonitor_37_or60;
  wire  TLMonitor_37_or29;
  wire  TLMonitor_37_or248;
  wire  TLMonitor_37_or123;
  wire  TLMonitor_37_or250;
  wire  TLMonitor_37_or124;
  wire  TLMonitor_37_or61;
  wire  TLMonitor_37_or252;
  wire  TLMonitor_37_or125;
  wire  TLMonitor_37_or254;
  wire  TLMonitor_37_or126;
  wire  TLMonitor_37_or62;
  wire  TLMonitor_37_or30;
  wire  TLMonitor_37_or14;
  wire  TLMonitor_37_or6;
  wire  TLMonitor_37_or2;
  wire  TLMonitor_37_or0;
  reg  TLMonitor_37_metaAssert;
  reg [31:0] _RAND_32;
  assign _T_4 = io_in_a_bits_source == 2'h0; // @[Parameters.scala 47:9]
  assign _T_5 = io_in_a_bits_source == 2'h1; // @[Parameters.scala 47:9]
  assign _T_6 = io_in_a_bits_source == 2'h2; // @[Parameters.scala 47:9]
  assign _T_8 = _T_4 | _T_5; // @[Parameters.scala 1016:46]
  assign _T_9 = _T_8 | _T_6; // @[Parameters.scala 1016:46]
  assign _T_11 = 27'hfff << io_in_a_bits_size; // @[package.scala 212:77]
  assign _GEN_71 = {{20'd0}, ~_T_11[11:0]}; // @[Edges.scala 22:16]
  assign _T_14 = io_in_a_bits_address & _GEN_71; // @[Edges.scala 22:16]
  assign _T_15 = _T_14 == 32'h0; // @[Edges.scala 22:24]
  assign _T_18 = 4'h1 << io_in_a_bits_size[1:0]; // @[OneHot.scala 65:12]
  assign _T_20 = _T_18[2:0] | 3'h1; // @[Misc.scala 201:81]
  assign _T_21 = io_in_a_bits_size >= 4'h3; // @[Misc.scala 205:21]
  assign _T_26 = _T_20[2] & ~io_in_a_bits_address[2]; // @[Misc.scala 214:38]
  assign _T_27 = _T_21 | _T_26; // @[Misc.scala 214:29]
  assign _T_29 = _T_20[2] & io_in_a_bits_address[2]; // @[Misc.scala 214:38]
  assign _T_30 = _T_21 | _T_29; // @[Misc.scala 214:29]
  assign _T_34 = ~io_in_a_bits_address[2] & ~io_in_a_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_35 = _T_20[1] & _T_34; // @[Misc.scala 214:38]
  assign _T_36 = _T_27 | _T_35; // @[Misc.scala 214:29]
  assign _T_37 = ~io_in_a_bits_address[2] & io_in_a_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_38 = _T_20[1] & _T_37; // @[Misc.scala 214:38]
  assign _T_39 = _T_27 | _T_38; // @[Misc.scala 214:29]
  assign _T_40 = io_in_a_bits_address[2] & ~io_in_a_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_41 = _T_20[1] & _T_40; // @[Misc.scala 214:38]
  assign _T_42 = _T_30 | _T_41; // @[Misc.scala 214:29]
  assign _T_43 = io_in_a_bits_address[2] & io_in_a_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_44 = _T_20[1] & _T_43; // @[Misc.scala 214:38]
  assign _T_45 = _T_30 | _T_44; // @[Misc.scala 214:29]
  assign _T_49 = _T_34 & ~io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_50 = _T_20[0] & _T_49; // @[Misc.scala 214:38]
  assign _T_51 = _T_36 | _T_50; // @[Misc.scala 214:29]
  assign _T_52 = _T_34 & io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_53 = _T_20[0] & _T_52; // @[Misc.scala 214:38]
  assign _T_54 = _T_36 | _T_53; // @[Misc.scala 214:29]
  assign _T_55 = _T_37 & ~io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_56 = _T_20[0] & _T_55; // @[Misc.scala 214:38]
  assign _T_57 = _T_39 | _T_56; // @[Misc.scala 214:29]
  assign _T_58 = _T_37 & io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_59 = _T_20[0] & _T_58; // @[Misc.scala 214:38]
  assign _T_60 = _T_39 | _T_59; // @[Misc.scala 214:29]
  assign _T_61 = _T_40 & ~io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_62 = _T_20[0] & _T_61; // @[Misc.scala 214:38]
  assign _T_63 = _T_42 | _T_62; // @[Misc.scala 214:29]
  assign _T_64 = _T_40 & io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_65 = _T_20[0] & _T_64; // @[Misc.scala 214:38]
  assign _T_66 = _T_42 | _T_65; // @[Misc.scala 214:29]
  assign _T_67 = _T_43 & ~io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_68 = _T_20[0] & _T_67; // @[Misc.scala 214:38]
  assign _T_69 = _T_45 | _T_68; // @[Misc.scala 214:29]
  assign _T_70 = _T_43 & io_in_a_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_71 = _T_20[0] & _T_70; // @[Misc.scala 214:38]
  assign _T_72 = _T_45 | _T_71; // @[Misc.scala 214:29]
  assign _T_79 = {_T_72,_T_69,_T_66,_T_63,_T_60,_T_57,_T_54,_T_51}; // @[Cat.scala 29:58]
  assign _T_83 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49]
  assign _T_109 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 82:25]
  assign _T_111 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 93:42]
  assign _T_118 = _T_111 & _T_9; // @[Parameters.scala 1066:30]
  assign _T_128 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 93:42]
  assign _T_131 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  assign _T_132 = {1'b0,$signed(_T_131)}; // @[Parameters.scala 137:49]
  assign _T_134 = $signed(_T_132) & 33'sh80000000; // @[Parameters.scala 137:52]
  assign _T_135 = $signed(_T_134) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_136 = _T_128 & _T_135; // @[Parameters.scala 601:56]
  assign _T_139 = _T_118 & _T_136; // @[Parameters.scala 1240:195]
  assign _T_141 = _T_139 | reset; // @[Monitor.scala 44:11]
  assign _T_147 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 92:48]
  assign _T_148 = _T_4 & _T_147; // @[Mux.scala 27:72]
  assign _T_165 = _T_148 & _T_111; // @[Parameters.scala 1255:195]
  assign _T_167 = _T_165 | reset; // @[Monitor.scala 44:11]
  assign _T_170 = _T_9 | reset; // @[Monitor.scala 44:11]
  assign _T_174 = _T_21 | reset; // @[Monitor.scala 44:11]
  assign _T_177 = _T_15 | reset; // @[Monitor.scala 44:11]
  assign _T_179 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 110:27]
  assign _T_181 = _T_179 | reset; // @[Monitor.scala 44:11]
  assign _T_184 = ~io_in_a_bits_mask == 8'h0; // @[Monitor.scala 89:31]
  assign _T_186 = _T_184 | reset; // @[Monitor.scala 44:11]
  assign _T_190 = ~io_in_a_bits_corrupt | reset; // @[Monitor.scala 44:11]
  assign _T_192 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 93:25]
  assign _T_266 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 100:31]
  assign _T_268 = _T_266 | reset; // @[Monitor.scala 44:11]
  assign _T_279 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 105:25]
  assign _T_294 = io_in_a_bits_address ^ 32'h2000; // @[Parameters.scala 137:31]
  assign _T_295 = {1'b0,$signed(_T_294)}; // @[Parameters.scala 137:49]
  assign _T_297 = $signed(_T_295) & 33'shca012000; // @[Parameters.scala 137:52]
  assign _T_298 = $signed(_T_297) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_299 = _T_111 & _T_298; // @[Parameters.scala 601:56]
  assign _T_307 = $signed(_T_83) & 33'shca012000; // @[Parameters.scala 137:52]
  assign _T_308 = $signed(_T_307) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_309 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31]
  assign _T_310 = {1'b0,$signed(_T_309)}; // @[Parameters.scala 137:49]
  assign _T_312 = $signed(_T_310) & 33'shca010000; // @[Parameters.scala 137:52]
  assign _T_313 = $signed(_T_312) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_314 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31]
  assign _T_315 = {1'b0,$signed(_T_314)}; // @[Parameters.scala 137:49]
  assign _T_317 = $signed(_T_315) & 33'shca010000; // @[Parameters.scala 137:52]
  assign _T_318 = $signed(_T_317) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_319 = io_in_a_bits_address ^ 32'h8000000; // @[Parameters.scala 137:31]
  assign _T_320 = {1'b0,$signed(_T_319)}; // @[Parameters.scala 137:49]
  assign _T_322 = $signed(_T_320) & 33'shc8000000; // @[Parameters.scala 137:52]
  assign _T_323 = $signed(_T_322) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_324 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  assign _T_325 = {1'b0,$signed(_T_324)}; // @[Parameters.scala 137:49]
  assign _T_327 = $signed(_T_325) & 33'shc0000000; // @[Parameters.scala 137:52]
  assign _T_328 = $signed(_T_327) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_332 = $signed(_T_132) & 33'shc0000000; // @[Parameters.scala 137:52]
  assign _T_333 = $signed(_T_332) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_334 = _T_308 | _T_313; // @[Parameters.scala 602:42]
  assign _T_335 = _T_334 | _T_318; // @[Parameters.scala 602:42]
  assign _T_336 = _T_335 | _T_323; // @[Parameters.scala 602:42]
  assign _T_337 = _T_336 | _T_328; // @[Parameters.scala 602:42]
  assign _T_338 = _T_337 | _T_333; // @[Parameters.scala 602:42]
  assign _T_339 = _T_128 & _T_338; // @[Parameters.scala 601:56]
  assign _T_341 = _T_299 | _T_339; // @[Parameters.scala 603:30]
  assign _T_342 = _T_118 & _T_341; // @[Parameters.scala 1243:195]
  assign _T_344 = _T_342 | reset; // @[Monitor.scala 44:11]
  assign _T_352 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31]
  assign _T_354 = _T_352 | reset; // @[Monitor.scala 44:11]
  assign _T_356 = io_in_a_bits_mask == _T_79; // @[Monitor.scala 110:30]
  assign _T_358 = _T_356 | reset; // @[Monitor.scala 44:11]
  assign _T_364 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  assign _T_409 = _T_308 | _T_318; // @[Parameters.scala 602:42]
  assign _T_410 = _T_409 | _T_323; // @[Parameters.scala 602:42]
  assign _T_411 = _T_410 | _T_333; // @[Parameters.scala 602:42]
  assign _T_412 = _T_128 & _T_411; // @[Parameters.scala 601:56]
  assign _T_421 = io_in_a_bits_size <= 4'h8; // @[Parameters.scala 93:42]
  assign _T_429 = _T_421 & _T_328; // @[Parameters.scala 601:56]
  assign _T_431 = _T_299 | _T_412; // @[Parameters.scala 603:30]
  assign _T_433 = _T_431 | _T_429; // @[Parameters.scala 603:30]
  assign _T_434 = _T_118 & _T_433; // @[Parameters.scala 1244:195]
  assign _T_436 = _T_434 | reset; // @[Monitor.scala 44:11]
  assign _T_452 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  assign _T_537 = io_in_a_bits_mask & ~_T_79; // @[Monitor.scala 127:31]
  assign _T_538 = _T_537 == 8'h0; // @[Monitor.scala 127:40]
  assign _T_540 = _T_538 | reset; // @[Monitor.scala 44:11]
  assign _T_542 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  assign _T_554 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 93:42]
  assign _T_560 = $signed(_T_83) & 33'shc8010000; // @[Parameters.scala 137:52]
  assign _T_561 = $signed(_T_560) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_567 = _T_561 | _T_323; // @[Parameters.scala 602:42]
  assign _T_568 = _T_554 & _T_567; // @[Parameters.scala 601:56]
  assign _T_590 = _T_118 & _T_568; // @[Parameters.scala 1241:195]
  assign _T_592 = _T_590 | reset; // @[Monitor.scala 44:11]
  assign _T_600 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 140:33]
  assign _T_602 = _T_600 | reset; // @[Monitor.scala 44:11]
  assign _T_608 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  assign _T_666 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 147:30]
  assign _T_668 = _T_666 | reset; // @[Monitor.scala 44:11]
  assign _T_674 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  assign _T_734 = _T_118 & _T_299; // @[Parameters.scala 1246:195]
  assign _T_736 = _T_734 | reset; // @[Monitor.scala 44:11]
  assign _T_744 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 160:28]
  assign _T_746 = _T_744 | reset; // @[Monitor.scala 44:11]
  assign _T_756 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 44:24]
  assign _T_758 = _T_756 | reset; // @[Monitor.scala 51:11]
  assign _T_760 = io_in_d_bits_source == 2'h0; // @[Parameters.scala 47:9]
  assign _T_761 = io_in_d_bits_source == 2'h1; // @[Parameters.scala 47:9]
  assign _T_762 = io_in_d_bits_source == 2'h2; // @[Parameters.scala 47:9]
  assign _T_764 = _T_760 | _T_761; // @[Parameters.scala 1016:46]
  assign _T_765 = _T_764 | _T_762; // @[Parameters.scala 1016:46]
  assign _T_767 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  assign _T_769 = _T_765 | reset; // @[Monitor.scala 51:11]
  assign _T_771 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27]
  assign _T_773 = _T_771 | reset; // @[Monitor.scala 51:11]
  assign _T_775 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  assign _T_777 = _T_775 | reset; // @[Monitor.scala 51:11]
  assign _T_781 = ~io_in_d_bits_corrupt | reset; // @[Monitor.scala 51:11]
  assign _T_785 = ~io_in_d_bits_denied | reset; // @[Monitor.scala 51:11]
  assign _T_787 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  assign _T_798 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 104:26]
  assign _T_800 = _T_798 | reset; // @[Monitor.scala 51:11]
  assign _T_802 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  assign _T_804 = _T_802 | reset; // @[Monitor.scala 51:11]
  assign _T_815 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  assign _T_835 = ~io_in_d_bits_denied | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  assign _T_837 = _T_835 | reset; // @[Monitor.scala 51:11]
  assign _T_844 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  assign _T_861 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  assign _T_879 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  assign _T_896 = io_in_b_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  assign _T_898 = _T_896 | reset; // @[Monitor.scala 44:11]
  assign _T_900 = io_in_b_bits_source == 2'h0; // @[Parameters.scala 47:9]
  assign _T_903 = {1'b0,$signed(io_in_b_bits_address)}; // @[Parameters.scala 137:49]
  assign _T_908 = io_in_b_bits_source == 2'h1; // @[Parameters.scala 47:9]
  assign _T_916 = io_in_b_bits_source == 2'h2; // @[Parameters.scala 47:9]
  assign _T_929 = io_in_b_bits_address ^ 32'h3000; // @[Parameters.scala 137:31]
  assign _T_930 = {1'b0,$signed(_T_929)}; // @[Parameters.scala 137:49]
  assign _T_932 = $signed(_T_930) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _T_933 = $signed(_T_932) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_934 = io_in_b_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31]
  assign _T_935 = {1'b0,$signed(_T_934)}; // @[Parameters.scala 137:49]
  assign _T_937 = $signed(_T_935) & -33'sh4000000; // @[Parameters.scala 137:52]
  assign _T_938 = $signed(_T_937) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_939 = io_in_b_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31]
  assign _T_940 = {1'b0,$signed(_T_939)}; // @[Parameters.scala 137:49]
  assign _T_942 = $signed(_T_940) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _T_943 = $signed(_T_942) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_947 = $signed(_T_903) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _T_948 = $signed(_T_947) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_949 = io_in_b_bits_address ^ 32'h10000; // @[Parameters.scala 137:31]
  assign _T_950 = {1'b0,$signed(_T_949)}; // @[Parameters.scala 137:49]
  assign _T_952 = $signed(_T_950) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _T_953 = $signed(_T_952) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_954 = io_in_b_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  assign _T_955 = {1'b0,$signed(_T_954)}; // @[Parameters.scala 137:49]
  assign _T_957 = $signed(_T_955) & -33'sh10000000; // @[Parameters.scala 137:52]
  assign _T_958 = $signed(_T_957) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_959 = io_in_b_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31]
  assign _T_960 = {1'b0,$signed(_T_959)}; // @[Parameters.scala 137:49]
  assign _T_962 = $signed(_T_960) & -33'sh20000000; // @[Parameters.scala 137:52]
  assign _T_963 = $signed(_T_962) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_965 = _T_933 | _T_938; // @[Parameters.scala 556:64]
  assign _T_966 = _T_965 | _T_943; // @[Parameters.scala 556:64]
  assign _T_967 = _T_966 | _T_948; // @[Parameters.scala 556:64]
  assign _T_968 = _T_967 | _T_953; // @[Parameters.scala 556:64]
  assign _T_969 = _T_968 | _T_958; // @[Parameters.scala 556:64]
  assign _T_970 = _T_969 | _T_963; // @[Parameters.scala 556:64]
  assign _T_972 = 27'hfff << io_in_b_bits_size; // @[package.scala 212:77]
  assign _GEN_72 = {{20'd0}, ~_T_972[11:0]}; // @[Edges.scala 22:16]
  assign _T_975 = io_in_b_bits_address & _GEN_72; // @[Edges.scala 22:16]
  assign _T_976 = _T_975 == 32'h0; // @[Edges.scala 22:24]
  assign _T_979 = 4'h1 << io_in_b_bits_size[1:0]; // @[OneHot.scala 65:12]
  assign _T_981 = _T_979[2:0] | 3'h1; // @[Misc.scala 201:81]
  assign _T_982 = io_in_b_bits_size >= 4'h3; // @[Misc.scala 205:21]
  assign _T_987 = _T_981[2] & ~io_in_b_bits_address[2]; // @[Misc.scala 214:38]
  assign _T_988 = _T_982 | _T_987; // @[Misc.scala 214:29]
  assign _T_990 = _T_981[2] & io_in_b_bits_address[2]; // @[Misc.scala 214:38]
  assign _T_991 = _T_982 | _T_990; // @[Misc.scala 214:29]
  assign _T_995 = ~io_in_b_bits_address[2] & ~io_in_b_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_996 = _T_981[1] & _T_995; // @[Misc.scala 214:38]
  assign _T_997 = _T_988 | _T_996; // @[Misc.scala 214:29]
  assign _T_998 = ~io_in_b_bits_address[2] & io_in_b_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_999 = _T_981[1] & _T_998; // @[Misc.scala 214:38]
  assign _T_1000 = _T_988 | _T_999; // @[Misc.scala 214:29]
  assign _T_1001 = io_in_b_bits_address[2] & ~io_in_b_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_1002 = _T_981[1] & _T_1001; // @[Misc.scala 214:38]
  assign _T_1003 = _T_991 | _T_1002; // @[Misc.scala 214:29]
  assign _T_1004 = io_in_b_bits_address[2] & io_in_b_bits_address[1]; // @[Misc.scala 213:27]
  assign _T_1005 = _T_981[1] & _T_1004; // @[Misc.scala 214:38]
  assign _T_1006 = _T_991 | _T_1005; // @[Misc.scala 214:29]
  assign _T_1010 = _T_995 & ~io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_1011 = _T_981[0] & _T_1010; // @[Misc.scala 214:38]
  assign _T_1012 = _T_997 | _T_1011; // @[Misc.scala 214:29]
  assign _T_1013 = _T_995 & io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_1014 = _T_981[0] & _T_1013; // @[Misc.scala 214:38]
  assign _T_1015 = _T_997 | _T_1014; // @[Misc.scala 214:29]
  assign _T_1016 = _T_998 & ~io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_1017 = _T_981[0] & _T_1016; // @[Misc.scala 214:38]
  assign _T_1018 = _T_1000 | _T_1017; // @[Misc.scala 214:29]
  assign _T_1019 = _T_998 & io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_1020 = _T_981[0] & _T_1019; // @[Misc.scala 214:38]
  assign _T_1021 = _T_1000 | _T_1020; // @[Misc.scala 214:29]
  assign _T_1022 = _T_1001 & ~io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_1023 = _T_981[0] & _T_1022; // @[Misc.scala 214:38]
  assign _T_1024 = _T_1003 | _T_1023; // @[Misc.scala 214:29]
  assign _T_1025 = _T_1001 & io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_1026 = _T_981[0] & _T_1025; // @[Misc.scala 214:38]
  assign _T_1027 = _T_1003 | _T_1026; // @[Misc.scala 214:29]
  assign _T_1028 = _T_1004 & ~io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_1029 = _T_981[0] & _T_1028; // @[Misc.scala 214:38]
  assign _T_1030 = _T_1006 | _T_1029; // @[Misc.scala 214:29]
  assign _T_1031 = _T_1004 & io_in_b_bits_address[0]; // @[Misc.scala 213:27]
  assign _T_1032 = _T_981[0] & _T_1031; // @[Misc.scala 214:38]
  assign _T_1033 = _T_1006 | _T_1032; // @[Misc.scala 214:29]
  assign _T_1040 = {_T_1033,_T_1030,_T_1027,_T_1024,_T_1021,_T_1018,_T_1015,_T_1012}; // @[Cat.scala 29:58]
  assign _T_1047 = _T_916 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  assign _GEN_73 = {{1'd0}, _T_908}; // @[Mux.scala 27:72]
  assign _T_1049 = _GEN_73 | _T_1047; // @[Mux.scala 27:72]
  assign _T_1051 = _T_1049 == io_in_b_bits_source; // @[Monitor.scala 165:113]
  assign _T_1052 = io_in_b_bits_opcode == 3'h6; // @[Monitor.scala 167:25]
  assign _T_1057 = 4'h6 == io_in_b_bits_size; // @[Parameters.scala 92:48]
  assign _T_1058 = _T_900 & _T_1057; // @[Mux.scala 27:72]
  assign _T_1065 = io_in_b_bits_size <= 4'hc; // @[Parameters.scala 93:42]
  assign _T_1075 = _T_1058 & _T_1065; // @[Parameters.scala 1255:195]
  assign _T_1077 = _T_1075 | reset; // @[Monitor.scala 44:11]
  assign _T_1080 = _T_970 | reset; // @[Monitor.scala 44:11]
  assign _T_1083 = _T_1051 | reset; // @[Monitor.scala 44:11]
  assign _T_1086 = _T_976 | reset; // @[Monitor.scala 44:11]
  assign _T_1088 = io_in_b_bits_param <= 2'h2; // @[Bundles.scala 104:26]
  assign _T_1090 = _T_1088 | reset; // @[Monitor.scala 44:11]
  assign _T_1092 = io_in_b_bits_mask == _T_1040; // @[Monitor.scala 173:30]
  assign _T_1094 = _T_1092 | reset; // @[Monitor.scala 44:11]
  assign _T_1098 = ~io_in_b_bits_corrupt | reset; // @[Monitor.scala 44:11]
  assign _T_1100 = io_in_b_bits_opcode == 3'h4; // @[Monitor.scala 177:25]
  assign _T_1125 = io_in_b_bits_param == 2'h0; // @[Monitor.scala 182:31]
  assign _T_1127 = _T_1125 | reset; // @[Monitor.scala 44:11]
  assign _T_1137 = io_in_b_bits_opcode == 3'h0; // @[Monitor.scala 187:25]
  assign _T_1170 = io_in_b_bits_opcode == 3'h1; // @[Monitor.scala 196:25]
  assign _T_1200 = io_in_b_bits_mask & ~_T_1040; // @[Monitor.scala 202:31]
  assign _T_1201 = _T_1200 == 8'h0; // @[Monitor.scala 202:40]
  assign _T_1203 = _T_1201 | reset; // @[Monitor.scala 44:11]
  assign _T_1205 = io_in_b_bits_opcode == 3'h2; // @[Monitor.scala 205:25]
  assign _T_1238 = io_in_b_bits_opcode == 3'h3; // @[Monitor.scala 214:25]
  assign _T_1271 = io_in_b_bits_opcode == 3'h5; // @[Monitor.scala 223:25]
  assign _T_1308 = io_in_c_bits_source == 2'h0; // @[Parameters.scala 47:9]
  assign _T_1309 = io_in_c_bits_source == 2'h1; // @[Parameters.scala 47:9]
  assign _T_1310 = io_in_c_bits_source == 2'h2; // @[Parameters.scala 47:9]
  assign _T_1312 = _T_1308 | _T_1309; // @[Parameters.scala 1016:46]
  assign _T_1313 = _T_1312 | _T_1310; // @[Parameters.scala 1016:46]
  assign _T_1315 = 27'hfff << io_in_c_bits_size; // @[package.scala 212:77]
  assign _GEN_74 = {{20'd0}, ~_T_1315[11:0]}; // @[Edges.scala 22:16]
  assign _T_1318 = io_in_c_bits_address & _GEN_74; // @[Edges.scala 22:16]
  assign _T_1319 = _T_1318 == 32'h0; // @[Edges.scala 22:24]
  assign _T_1320 = io_in_c_bits_address ^ 32'h3000; // @[Parameters.scala 137:31]
  assign _T_1321 = {1'b0,$signed(_T_1320)}; // @[Parameters.scala 137:49]
  assign _T_1323 = $signed(_T_1321) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _T_1324 = $signed(_T_1323) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1325 = io_in_c_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31]
  assign _T_1326 = {1'b0,$signed(_T_1325)}; // @[Parameters.scala 137:49]
  assign _T_1328 = $signed(_T_1326) & -33'sh4000000; // @[Parameters.scala 137:52]
  assign _T_1329 = $signed(_T_1328) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1330 = io_in_c_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31]
  assign _T_1331 = {1'b0,$signed(_T_1330)}; // @[Parameters.scala 137:49]
  assign _T_1333 = $signed(_T_1331) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _T_1334 = $signed(_T_1333) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1336 = {1'b0,$signed(io_in_c_bits_address)}; // @[Parameters.scala 137:49]
  assign _T_1338 = $signed(_T_1336) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _T_1339 = $signed(_T_1338) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1340 = io_in_c_bits_address ^ 32'h10000; // @[Parameters.scala 137:31]
  assign _T_1341 = {1'b0,$signed(_T_1340)}; // @[Parameters.scala 137:49]
  assign _T_1343 = $signed(_T_1341) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _T_1344 = $signed(_T_1343) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1345 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  assign _T_1346 = {1'b0,$signed(_T_1345)}; // @[Parameters.scala 137:49]
  assign _T_1348 = $signed(_T_1346) & -33'sh10000000; // @[Parameters.scala 137:52]
  assign _T_1349 = $signed(_T_1348) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1350 = io_in_c_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31]
  assign _T_1351 = {1'b0,$signed(_T_1350)}; // @[Parameters.scala 137:49]
  assign _T_1353 = $signed(_T_1351) & -33'sh20000000; // @[Parameters.scala 137:52]
  assign _T_1354 = $signed(_T_1353) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1356 = _T_1324 | _T_1329; // @[Parameters.scala 556:64]
  assign _T_1357 = _T_1356 | _T_1334; // @[Parameters.scala 556:64]
  assign _T_1358 = _T_1357 | _T_1339; // @[Parameters.scala 556:64]
  assign _T_1359 = _T_1358 | _T_1344; // @[Parameters.scala 556:64]
  assign _T_1360 = _T_1359 | _T_1349; // @[Parameters.scala 556:64]
  assign _T_1361 = _T_1360 | _T_1354; // @[Parameters.scala 556:64]
  assign _T_1391 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 242:25]
  assign _T_1393 = _T_1361 | reset; // @[Monitor.scala 44:11]
  assign _T_1396 = _T_1313 | reset; // @[Monitor.scala 44:11]
  assign _T_1398 = io_in_c_bits_size >= 4'h3; // @[Monitor.scala 245:30]
  assign _T_1400 = _T_1398 | reset; // @[Monitor.scala 44:11]
  assign _T_1403 = _T_1319 | reset; // @[Monitor.scala 44:11]
  assign _T_1405 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 122:29]
  assign _T_1407 = _T_1405 | reset; // @[Monitor.scala 44:11]
  assign _T_1413 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 251:25]
  assign _T_1431 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 259:25]
  assign _T_1433 = io_in_c_bits_size <= 4'hc; // @[Parameters.scala 93:42]
  assign _T_1440 = _T_1433 & _T_1313; // @[Parameters.scala 1066:30]
  assign _T_1450 = io_in_c_bits_size <= 4'h6; // @[Parameters.scala 93:42]
  assign _T_1456 = $signed(_T_1346) & 33'sh80000000; // @[Parameters.scala 137:52]
  assign _T_1457 = $signed(_T_1456) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_1458 = _T_1450 & _T_1457; // @[Parameters.scala 601:56]
  assign _T_1461 = _T_1440 & _T_1458; // @[Parameters.scala 1240:195]
  assign _T_1463 = _T_1461 | reset; // @[Monitor.scala 44:11]
  assign _T_1469 = 4'h6 == io_in_c_bits_size; // @[Parameters.scala 92:48]
  assign _T_1470 = _T_1308 & _T_1469; // @[Mux.scala 27:72]
  assign _T_1487 = _T_1470 & _T_1433; // @[Parameters.scala 1255:195]
  assign _T_1489 = _T_1487 | reset; // @[Monitor.scala 44:11]
  assign _T_1501 = io_in_c_bits_param <= 3'h2; // @[Bundles.scala 116:29]
  assign _T_1503 = _T_1501 | reset; // @[Monitor.scala 44:11]
  assign _T_1509 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 269:25]
  assign _T_1583 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 278:25]
  assign _T_1593 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 282:31]
  assign _T_1595 = _T_1593 | reset; // @[Monitor.scala 44:11]
  assign _T_1601 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 286:25]
  assign _T_1615 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 293:25]
  assign _T_1637 = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  assign _T_1642 = ~_T_11[11:3]; // @[Edges.scala 221:59]
  assign _T_1648 = _T_1646 - 9'h1; // @[Edges.scala 231:28]
  assign _T_1649 = _T_1646 == 9'h0; // @[Edges.scala 232:25]
  assign _T_1663 = io_in_a_valid & ~_T_1649; // @[Monitor.scala 389:19]
  assign _T_1664 = io_in_a_bits_opcode == _T_1657; // @[Monitor.scala 390:32]
  assign _T_1666 = _T_1664 | reset; // @[Monitor.scala 44:11]
  assign _T_1668 = io_in_a_bits_param == _T_1658; // @[Monitor.scala 391:32]
  assign _T_1670 = _T_1668 | reset; // @[Monitor.scala 44:11]
  assign _T_1672 = io_in_a_bits_size == _T_1659; // @[Monitor.scala 392:32]
  assign _T_1674 = _T_1672 | reset; // @[Monitor.scala 44:11]
  assign _T_1676 = io_in_a_bits_source == _T_1660; // @[Monitor.scala 393:32]
  assign _T_1678 = _T_1676 | reset; // @[Monitor.scala 44:11]
  assign _T_1680 = io_in_a_bits_address == _T_1661; // @[Monitor.scala 394:32]
  assign _T_1682 = _T_1680 | reset; // @[Monitor.scala 44:11]
  assign _T_1685 = _T_1637 & _T_1649; // @[Monitor.scala 396:20]
  assign _T_1686 = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  assign _T_1688 = 27'hfff << io_in_d_bits_size; // @[package.scala 212:77]
  assign _T_1691 = ~_T_1688[11:3]; // @[Edges.scala 221:59]
  assign _T_1696 = _T_1694 - 9'h1; // @[Edges.scala 231:28]
  assign _T_1697 = _T_1694 == 9'h0; // @[Edges.scala 232:25]
  assign _T_1712 = io_in_d_valid & ~_T_1697; // @[Monitor.scala 541:19]
  assign _T_1713 = io_in_d_bits_opcode == _T_1705; // @[Monitor.scala 542:29]
  assign _T_1715 = _T_1713 | reset; // @[Monitor.scala 51:11]
  assign _T_1717 = io_in_d_bits_param == _T_1706; // @[Monitor.scala 543:29]
  assign _T_1719 = _T_1717 | reset; // @[Monitor.scala 51:11]
  assign _T_1721 = io_in_d_bits_size == _T_1707; // @[Monitor.scala 544:29]
  assign _T_1723 = _T_1721 | reset; // @[Monitor.scala 51:11]
  assign _T_1725 = io_in_d_bits_source == _T_1708; // @[Monitor.scala 545:29]
  assign _T_1727 = _T_1725 | reset; // @[Monitor.scala 51:11]
  assign _T_1729 = io_in_d_bits_sink == _T_1709; // @[Monitor.scala 546:29]
  assign _T_1731 = _T_1729 | reset; // @[Monitor.scala 51:11]
  assign _T_1733 = io_in_d_bits_denied == _T_1710; // @[Monitor.scala 547:29]
  assign _T_1735 = _T_1733 | reset; // @[Monitor.scala 51:11]
  assign _T_1738 = _T_1686 & _T_1697; // @[Monitor.scala 549:20]
  assign _T_1739 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37]
  assign _T_1750 = _T_1748 - 9'h1; // @[Edges.scala 231:28]
  assign _T_1751 = _T_1748 == 9'h0; // @[Edges.scala 232:25]
  assign _T_1765 = io_in_b_valid & ~_T_1751; // @[Monitor.scala 412:19]
  assign _T_1766 = io_in_b_bits_opcode == _T_1759; // @[Monitor.scala 413:32]
  assign _T_1768 = _T_1766 | reset; // @[Monitor.scala 44:11]
  assign _T_1770 = io_in_b_bits_param == _T_1760; // @[Monitor.scala 414:32]
  assign _T_1772 = _T_1770 | reset; // @[Monitor.scala 44:11]
  assign _T_1774 = io_in_b_bits_size == _T_1761; // @[Monitor.scala 415:32]
  assign _T_1776 = _T_1774 | reset; // @[Monitor.scala 44:11]
  assign _T_1778 = io_in_b_bits_source == _T_1762; // @[Monitor.scala 416:32]
  assign _T_1780 = _T_1778 | reset; // @[Monitor.scala 44:11]
  assign _T_1782 = io_in_b_bits_address == _T_1763; // @[Monitor.scala 417:32]
  assign _T_1784 = _T_1782 | reset; // @[Monitor.scala 44:11]
  assign _T_1787 = _T_1739 & _T_1751; // @[Monitor.scala 419:20]
  assign _T_1788 = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37]
  assign _T_1793 = ~_T_1315[11:3]; // @[Edges.scala 221:59]
  assign _T_1798 = _T_1796 - 9'h1; // @[Edges.scala 231:28]
  assign _T_1799 = _T_1796 == 9'h0; // @[Edges.scala 232:25]
  assign _T_1813 = io_in_c_valid & ~_T_1799; // @[Monitor.scala 517:19]
  assign _T_1814 = io_in_c_bits_opcode == _T_1807; // @[Monitor.scala 518:32]
  assign _T_1816 = _T_1814 | reset; // @[Monitor.scala 44:11]
  assign _T_1818 = io_in_c_bits_param == _T_1808; // @[Monitor.scala 519:32]
  assign _T_1820 = _T_1818 | reset; // @[Monitor.scala 44:11]
  assign _T_1822 = io_in_c_bits_size == _T_1809; // @[Monitor.scala 520:32]
  assign _T_1824 = _T_1822 | reset; // @[Monitor.scala 44:11]
  assign _T_1826 = io_in_c_bits_source == _T_1810; // @[Monitor.scala 521:32]
  assign _T_1828 = _T_1826 | reset; // @[Monitor.scala 44:11]
  assign _T_1830 = io_in_c_bits_address == _T_1811; // @[Monitor.scala 522:32]
  assign _T_1832 = _T_1830 | reset; // @[Monitor.scala 44:11]
  assign _T_1835 = _T_1788 & _T_1799; // @[Monitor.scala 524:20]
  assign _T_1847 = _T_1845 - 9'h1; // @[Edges.scala 231:28]
  assign a_first = _T_1845 == 9'h0; // @[Edges.scala 232:25]
  assign _T_1865 = _T_1863 - 9'h1; // @[Edges.scala 231:28]
  assign d_first = _T_1863 == 9'h0; // @[Edges.scala 232:25]
  assign _GEN_75 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 632:69]
  assign _T_1873 = {{1'd0}, _GEN_75}; // @[Monitor.scala 632:69]
  assign _T_1874 = inflight_opcodes >> _T_1873; // @[Monitor.scala 632:44]
  assign _T_1878 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  assign _GEN_76 = {{4'd0}, _T_1874}; // @[Monitor.scala 632:97]
  assign _T_1879 = _GEN_76 & _T_1878; // @[Monitor.scala 632:97]
  assign _T_1880 = {{1'd0}, _T_1879[15:1]}; // @[Monitor.scala 632:152]
  assign _T_1881 = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 636:65]
  assign _T_1882 = inflight_sizes >> _T_1881; // @[Monitor.scala 636:40]
  assign _T_1886 = 16'h100 - 16'h1; // @[Monitor.scala 609:57]
  assign _GEN_78 = {{8'd0}, _T_1886}; // @[Monitor.scala 636:91]
  assign _T_1887 = _T_1882 & _GEN_78; // @[Monitor.scala 636:91]
  assign _T_1888 = {{1'd0}, _T_1887[23:1]}; // @[Monitor.scala 636:144]
  assign _T_1892 = _T_1637 & a_first; // @[Monitor.scala 646:27]
  assign _T_1894 = 4'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  assign _T_1895 = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 648:53]
  assign _T_1896 = _T_1895 | 4'h1; // @[Monitor.scala 648:61]
  assign _T_1897 = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 649:49]
  assign _T_1898 = _T_1897 | 5'h1; // @[Monitor.scala 649:57]
  assign _GEN_80 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 650:72]
  assign _T_1899 = {{1'd0}, _GEN_80}; // @[Monitor.scala 650:72]
  assign a_opcodes_set_interm = _T_1892 ? _T_1896 : 4'h0; // @[Monitor.scala 646:72]
  assign _GEN_81 = {{31'd0}, a_opcodes_set_interm}; // @[Monitor.scala 650:47]
  assign _T_1900 = _GEN_81 << _T_1899; // @[Monitor.scala 650:47]
  assign _T_1901 = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 651:68]
  assign a_sizes_set_interm = _T_1892 ? _T_1898 : 5'h0; // @[Monitor.scala 646:72]
  assign _GEN_82 = {{31'd0}, a_sizes_set_interm}; // @[Monitor.scala 651:43]
  assign _T_1902 = _GEN_82 << _T_1901; // @[Monitor.scala 651:43]
  assign _T_1903 = inflight >> io_in_a_bits_source; // @[Monitor.scala 652:26]
  assign _T_1907 = ~_T_1903[0] | reset; // @[Monitor.scala 44:11]
  assign _GEN_27 = _T_1892 ? _T_1894 : 4'h0; // @[Monitor.scala 646:72]
  assign _GEN_30 = _T_1892 ? _T_1900 : 35'h0; // @[Monitor.scala 646:72]
  assign _GEN_31 = _T_1892 ? _T_1902 : 36'h0; // @[Monitor.scala 646:72]
  assign _T_1911 = _T_1686 & d_first; // @[Monitor.scala 663:27]
  assign _T_1914 = _T_1911 & ~_T_767; // @[Monitor.scala 663:72]
  assign _T_1915 = 4'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  assign _GEN_84 = {{31'd0}, _T_1878}; // @[Monitor.scala 665:76]
  assign _T_1921 = _GEN_84 << _T_1873; // @[Monitor.scala 665:76]
  assign _GEN_85 = {{31'd0}, _T_1886}; // @[Monitor.scala 666:72]
  assign _T_1927 = _GEN_85 << _T_1881; // @[Monitor.scala 666:72]
  assign _GEN_32 = _T_1914 ? _T_1915 : 4'h0; // @[Monitor.scala 663:91]
  assign _GEN_33 = _T_1914 ? _T_1921 : 47'h0; // @[Monitor.scala 663:91]
  assign _GEN_34 = _T_1914 ? _T_1927 : 47'h0; // @[Monitor.scala 663:91]
  assign _T_1928 = io_in_d_valid & d_first; // @[Monitor.scala 668:26]
  assign _T_1931 = _T_1928 & ~_T_767; // @[Monitor.scala 668:71]
  assign _T_1932 = inflight >> io_in_d_bits_source; // @[Monitor.scala 669:25]
  assign _T_1934 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 669:93]
  assign _T_1935 = io_in_a_valid & _T_1934; // @[Monitor.scala 669:68]
  assign _T_1936 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 669:142]
  assign _T_1937 = _T_1935 & _T_1936; // @[Monitor.scala 669:119]
  assign _T_1938 = _T_1937 & a_first; // @[Monitor.scala 669:166]
  assign _T_1939 = _T_1932[0] | _T_1938; // @[Monitor.scala 669:49]
  assign _T_1941 = _T_1939 | reset; // @[Monitor.scala 51:11]
  assign a_opcode_lookup = _T_1880[3:0]; // @[Monitor.scala 632:21]
  assign _GEN_37 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 670:37]
  assign _GEN_38 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_37; // @[Monitor.scala 670:37]
  assign _GEN_39 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_38; // @[Monitor.scala 670:37]
  assign _GEN_40 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_39; // @[Monitor.scala 670:37]
  assign _GEN_41 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_40; // @[Monitor.scala 670:37]
  assign _GEN_42 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_41; // @[Monitor.scala 670:37]
  assign _T_1944 = io_in_d_bits_opcode == _GEN_42; // @[Monitor.scala 670:37]
  assign _GEN_49 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_40; // @[Monitor.scala 670:96]
  assign _GEN_50 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_49; // @[Monitor.scala 670:96]
  assign _T_1946 = io_in_d_bits_opcode == _GEN_50; // @[Monitor.scala 670:96]
  assign _T_1947 = _T_1944 | _T_1946; // @[Monitor.scala 670:71]
  assign _GEN_53 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 671:60]
  assign _GEN_54 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_53; // @[Monitor.scala 671:60]
  assign _GEN_55 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_54; // @[Monitor.scala 671:60]
  assign _GEN_56 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_55; // @[Monitor.scala 671:60]
  assign _GEN_57 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_56; // @[Monitor.scala 671:60]
  assign _GEN_58 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_57; // @[Monitor.scala 671:60]
  assign _T_1948 = io_in_d_bits_opcode == _GEN_58; // @[Monitor.scala 671:60]
  assign _GEN_65 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_56; // @[Monitor.scala 671:124]
  assign _GEN_66 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_65; // @[Monitor.scala 671:124]
  assign _T_1949 = io_in_d_bits_opcode == _GEN_66; // @[Monitor.scala 671:124]
  assign _T_1950 = _T_1948 | _T_1949; // @[Monitor.scala 671:99]
  assign _T_1951 = io_in_a_valid & _T_1950; // @[Monitor.scala 671:34]
  assign _T_1952 = _T_1947 | _T_1951; // @[Monitor.scala 671:15]
  assign _T_1954 = _T_1952 | reset; // @[Monitor.scala 51:11]
  assign a_size_lookup = _T_1888[7:0]; // @[Monitor.scala 636:19]
  assign _GEN_86 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 673:34]
  assign _T_1956 = _GEN_86 == a_size_lookup; // @[Monitor.scala 673:34]
  assign _T_1958 = io_in_a_valid & _T_1936; // @[Monitor.scala 673:72]
  assign _T_1959 = _T_1956 | _T_1958; // @[Monitor.scala 673:53]
  assign _T_1961 = _T_1959 | reset; // @[Monitor.scala 51:11]
  assign _T_1964 = _T_1928 & a_first; // @[Monitor.scala 675:36]
  assign _T_1965 = _T_1964 & io_in_a_valid; // @[Monitor.scala 675:47]
  assign _T_1967 = _T_1965 & _T_1934; // @[Monitor.scala 675:65]
  assign _T_1969 = _T_1967 & ~_T_767; // @[Monitor.scala 675:116]
  assign _T_1971 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 676:32]
  assign _T_1973 = _T_1971 | reset; // @[Monitor.scala 51:11]
  assign a_set = _GEN_27[2:0]; // @[Monitor.scala 647:13]
  assign d_clr = _GEN_32[2:0]; // @[Monitor.scala 664:13]
  assign _T_1975 = a_set != d_clr; // @[Monitor.scala 680:20]
  assign _T_1976 = |a_set; // @[Monitor.scala 680:40]
  assign _T_1978 = _T_1975 | ~_T_1976; // @[Monitor.scala 680:30]
  assign _T_1980 = _T_1978 | reset; // @[Monitor.scala 51:11]
  assign _T_1982 = inflight | a_set; // @[Monitor.scala 683:27]
  assign _T_1984 = _T_1982 & ~d_clr; // @[Monitor.scala 683:36]
  assign a_opcodes_set = _GEN_30[11:0]; // @[Monitor.scala 650:21]
  assign _T_1985 = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 684:43]
  assign d_opcodes_clr = _GEN_33[11:0]; // @[Monitor.scala 665:21]
  assign _T_1987 = _T_1985 & ~d_opcodes_clr; // @[Monitor.scala 684:60]
  assign a_sizes_set = _GEN_31[23:0]; // @[Monitor.scala 651:19]
  assign _T_1988 = inflight_sizes | a_sizes_set; // @[Monitor.scala 685:39]
  assign d_sizes_clr = _GEN_34[23:0]; // @[Monitor.scala 666:19]
  assign _T_1990 = _T_1988 & ~d_sizes_clr; // @[Monitor.scala 685:54]
  assign _T_2017 = _T_2015 - 9'h1; // @[Edges.scala 231:28]
  assign _T_2018 = _T_2015 == 9'h0; // @[Edges.scala 232:25]
  assign _T_2028 = _T_1686 & _T_2018; // @[Monitor.scala 703:27]
  assign _T_2032 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 72:40]
  assign _T_2033 = _T_2028 & _T_2032; // @[Monitor.scala 703:38]
  assign _T_2034 = 4'h1 << io_in_d_bits_sink; // @[OneHot.scala 58:35]
  assign _T_2035 = _T_2006 >> io_in_d_bits_sink; // @[Monitor.scala 705:23]
  assign _T_2039 = ~_T_2035[0] | reset; // @[Monitor.scala 51:11]
  assign _GEN_69 = _T_2033 ? _T_2034 : 4'h0; // @[Monitor.scala 703:72]
  assign _T_2042 = io_in_e_ready & io_in_e_valid; // @[Decoupled.scala 40:37]
  assign _T_2045 = 4'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35]
  assign _T_2046 = _GEN_69 | _T_2006; // @[Monitor.scala 711:24]
  assign _T_2047 = _T_2046 >> io_in_e_bits_sink; // @[Monitor.scala 711:35]
  assign _T_2050 = _T_2047[0] | reset; // @[Monitor.scala 44:11]
  assign _GEN_70 = _T_2042 ? _T_2045 : 4'h0; // @[Monitor.scala 709:73]
  assign _T_2052 = _T_2006 | _GEN_69; // @[Monitor.scala 716:27]
  assign _T_2054 = _T_2052 & ~_GEN_70; // @[Monitor.scala 716:36]
  assign _GEN_87 = io_in_a_valid & _T_109; // @[Monitor.scala 44:11]
  assign _GEN_103 = io_in_a_valid & _T_192; // @[Monitor.scala 44:11]
  assign _GEN_121 = io_in_a_valid & _T_279; // @[Monitor.scala 44:11]
  assign _GEN_133 = io_in_a_valid & _T_364; // @[Monitor.scala 44:11]
  assign _GEN_143 = io_in_a_valid & _T_452; // @[Monitor.scala 44:11]
  assign _GEN_153 = io_in_a_valid & _T_542; // @[Monitor.scala 44:11]
  assign _GEN_163 = io_in_a_valid & _T_608; // @[Monitor.scala 44:11]
  assign _GEN_173 = io_in_a_valid & _T_674; // @[Monitor.scala 44:11]
  assign _GEN_185 = io_in_d_valid & _T_767; // @[Monitor.scala 51:11]
  assign _GEN_195 = io_in_d_valid & _T_787; // @[Monitor.scala 51:11]
  assign _GEN_205 = io_in_d_valid & _T_815; // @[Monitor.scala 51:11]
  assign _GEN_215 = io_in_d_valid & _T_844; // @[Monitor.scala 51:11]
  assign _GEN_221 = io_in_d_valid & _T_861; // @[Monitor.scala 51:11]
  assign _GEN_227 = io_in_d_valid & _T_879; // @[Monitor.scala 51:11]
  assign _GEN_233 = io_in_b_valid & _T_1052; // @[Monitor.scala 44:11]
  assign _GEN_247 = io_in_b_valid & _T_1100; // @[Monitor.scala 44:11]
  assign _GEN_261 = io_in_b_valid & _T_1137; // @[Monitor.scala 44:11]
  assign _GEN_273 = io_in_b_valid & _T_1170; // @[Monitor.scala 44:11]
  assign _GEN_285 = io_in_b_valid & _T_1205; // @[Monitor.scala 44:11]
  assign _GEN_295 = io_in_b_valid & _T_1238; // @[Monitor.scala 44:11]
  assign _GEN_305 = io_in_b_valid & _T_1271; // @[Monitor.scala 44:11]
  assign _GEN_317 = io_in_c_valid & _T_1391; // @[Monitor.scala 44:11]
  assign _GEN_327 = io_in_c_valid & _T_1413; // @[Monitor.scala 44:11]
  assign _GEN_337 = io_in_c_valid & _T_1431; // @[Monitor.scala 44:11]
  assign _GEN_349 = io_in_c_valid & _T_1509; // @[Monitor.scala 44:11]
  assign _GEN_361 = io_in_c_valid & _T_1583; // @[Monitor.scala 44:11]
  assign _GEN_369 = io_in_c_valid & _T_1601; // @[Monitor.scala 44:11]
  assign _GEN_377 = io_in_c_valid & _T_1615; // @[Monitor.scala 44:11]
  assign TLMonitor_37_covSum = 30'h0;
  assign io_covSum = TLMonitor_37_covSum;
  assign stopEn0 = _GEN_87 & ~_T_141;
  assign stopEn1 = _GEN_87 & ~_T_167;
  assign stopEn2 = _GEN_87 & ~_T_170;
  assign stopEn3 = _GEN_87 & ~_T_174;
  assign stopEn4 = _GEN_87 & ~_T_177;
  assign stopEn5 = _GEN_87 & ~_T_181;
  assign stopEn6 = _GEN_87 & ~_T_186;
  assign stopEn7 = _GEN_87 & ~_T_190;
  assign stopEn8 = _GEN_103 & ~_T_141;
  assign stopEn9 = _GEN_103 & ~_T_167;
  assign stopEn10 = _GEN_103 & ~_T_170;
  assign stopEn11 = _GEN_103 & ~_T_174;
  assign stopEn12 = _GEN_103 & ~_T_177;
  assign stopEn13 = _GEN_103 & ~_T_181;
  assign stopEn14 = _GEN_103 & ~_T_268;
  assign stopEn15 = _GEN_103 & ~_T_186;
  assign stopEn16 = _GEN_103 & ~_T_190;
  assign stopEn17 = _GEN_121 & ~_T_344;
  assign stopEn18 = _GEN_121 & ~_T_170;
  assign stopEn19 = _GEN_121 & ~_T_177;
  assign stopEn20 = _GEN_121 & ~_T_354;
  assign stopEn21 = _GEN_121 & ~_T_358;
  assign stopEn22 = _GEN_121 & ~_T_190;
  assign stopEn23 = _GEN_133 & ~_T_436;
  assign stopEn24 = _GEN_133 & ~_T_170;
  assign stopEn25 = _GEN_133 & ~_T_177;
  assign stopEn26 = _GEN_133 & ~_T_354;
  assign stopEn27 = _GEN_133 & ~_T_358;
  assign stopEn28 = _GEN_143 & ~_T_436;
  assign stopEn29 = _GEN_143 & ~_T_170;
  assign stopEn30 = _GEN_143 & ~_T_177;
  assign stopEn31 = _GEN_143 & ~_T_354;
  assign stopEn32 = _GEN_143 & ~_T_540;
  assign stopEn33 = _GEN_153 & ~_T_592;
  assign stopEn34 = _GEN_153 & ~_T_170;
  assign stopEn35 = _GEN_153 & ~_T_177;
  assign stopEn36 = _GEN_153 & ~_T_602;
  assign stopEn37 = _GEN_153 & ~_T_358;
  assign stopEn38 = _GEN_163 & ~_T_592;
  assign stopEn39 = _GEN_163 & ~_T_170;
  assign stopEn40 = _GEN_163 & ~_T_177;
  assign stopEn41 = _GEN_163 & ~_T_668;
  assign stopEn42 = _GEN_163 & ~_T_358;
  assign stopEn43 = _GEN_173 & ~_T_736;
  assign stopEn44 = _GEN_173 & ~_T_170;
  assign stopEn45 = _GEN_173 & ~_T_177;
  assign stopEn46 = _GEN_173 & ~_T_746;
  assign stopEn47 = _GEN_173 & ~_T_358;
  assign stopEn48 = _GEN_173 & ~_T_190;
  assign stopEn49 = io_in_d_valid & ~_T_758;
  assign stopEn50 = _GEN_185 & ~_T_769;
  assign stopEn51 = _GEN_185 & ~_T_773;
  assign stopEn52 = _GEN_185 & ~_T_777;
  assign stopEn53 = _GEN_185 & ~_T_781;
  assign stopEn54 = _GEN_185 & ~_T_785;
  assign stopEn55 = _GEN_195 & ~_T_769;
  assign stopEn56 = _GEN_195 & ~_T_773;
  assign stopEn57 = _GEN_195 & ~_T_800;
  assign stopEn58 = _GEN_195 & ~_T_804;
  assign stopEn59 = _GEN_195 & ~_T_781;
  assign stopEn60 = _GEN_205 & ~_T_769;
  assign stopEn61 = _GEN_205 & ~_T_773;
  assign stopEn62 = _GEN_205 & ~_T_800;
  assign stopEn63 = _GEN_205 & ~_T_804;
  assign stopEn64 = _GEN_205 & ~_T_837;
  assign stopEn65 = _GEN_215 & ~_T_769;
  assign stopEn66 = _GEN_215 & ~_T_777;
  assign stopEn67 = _GEN_215 & ~_T_781;
  assign stopEn68 = _GEN_221 & ~_T_769;
  assign stopEn69 = _GEN_221 & ~_T_777;
  assign stopEn70 = _GEN_221 & ~_T_837;
  assign stopEn71 = _GEN_227 & ~_T_769;
  assign stopEn72 = _GEN_227 & ~_T_777;
  assign stopEn73 = _GEN_227 & ~_T_781;
  assign stopEn74 = io_in_b_valid & ~_T_898;
  assign stopEn75 = _GEN_233 & ~_T_1077;
  assign stopEn76 = _GEN_233 & ~_T_1080;
  assign stopEn77 = _GEN_233 & ~_T_1083;
  assign stopEn78 = _GEN_233 & ~_T_1086;
  assign stopEn79 = _GEN_233 & ~_T_1090;
  assign stopEn80 = _GEN_233 & ~_T_1094;
  assign stopEn81 = _GEN_233 & ~_T_1098;
  assign stopEn82 = _GEN_247 & ~reset;
  assign stopEn83 = _GEN_247 & ~_T_1080;
  assign stopEn84 = _GEN_247 & ~_T_1083;
  assign stopEn85 = _GEN_247 & ~_T_1086;
  assign stopEn86 = _GEN_247 & ~_T_1127;
  assign stopEn87 = _GEN_247 & ~_T_1094;
  assign stopEn88 = _GEN_247 & ~_T_1098;
  assign stopEn89 = _GEN_261 & ~reset;
  assign stopEn90 = _GEN_261 & ~_T_1080;
  assign stopEn91 = _GEN_261 & ~_T_1083;
  assign stopEn92 = _GEN_261 & ~_T_1086;
  assign stopEn93 = _GEN_261 & ~_T_1127;
  assign stopEn94 = _GEN_261 & ~_T_1094;
  assign stopEn95 = _GEN_273 & ~reset;
  assign stopEn96 = _GEN_273 & ~_T_1080;
  assign stopEn97 = _GEN_273 & ~_T_1083;
  assign stopEn98 = _GEN_273 & ~_T_1086;
  assign stopEn99 = _GEN_273 & ~_T_1127;
  assign stopEn100 = _GEN_273 & ~_T_1203;
  assign stopEn101 = _GEN_285 & ~reset;
  assign stopEn102 = _GEN_285 & ~_T_1080;
  assign stopEn103 = _GEN_285 & ~_T_1083;
  assign stopEn104 = _GEN_285 & ~_T_1086;
  assign stopEn105 = _GEN_285 & ~_T_1094;
  assign stopEn106 = _GEN_295 & ~reset;
  assign stopEn107 = _GEN_295 & ~_T_1080;
  assign stopEn108 = _GEN_295 & ~_T_1083;
  assign stopEn109 = _GEN_295 & ~_T_1086;
  assign stopEn110 = _GEN_295 & ~_T_1094;
  assign stopEn111 = _GEN_305 & ~reset;
  assign stopEn112 = _GEN_305 & ~_T_1080;
  assign stopEn113 = _GEN_305 & ~_T_1083;
  assign stopEn114 = _GEN_305 & ~_T_1086;
  assign stopEn115 = _GEN_305 & ~_T_1094;
  assign stopEn116 = _GEN_305 & ~_T_1098;
  assign stopEn117 = _GEN_317 & ~_T_1393;
  assign stopEn118 = _GEN_317 & ~_T_1396;
  assign stopEn119 = _GEN_317 & ~_T_1400;
  assign stopEn120 = _GEN_317 & ~_T_1403;
  assign stopEn121 = _GEN_317 & ~_T_1407;
  assign stopEn122 = _GEN_327 & ~_T_1393;
  assign stopEn123 = _GEN_327 & ~_T_1396;
  assign stopEn124 = _GEN_327 & ~_T_1400;
  assign stopEn125 = _GEN_327 & ~_T_1403;
  assign stopEn126 = _GEN_327 & ~_T_1407;
  assign stopEn127 = _GEN_337 & ~_T_1463;
  assign stopEn128 = _GEN_337 & ~_T_1489;
  assign stopEn129 = _GEN_337 & ~_T_1396;
  assign stopEn130 = _GEN_337 & ~_T_1400;
  assign stopEn131 = _GEN_337 & ~_T_1403;
  assign stopEn132 = _GEN_337 & ~_T_1503;
  assign stopEn133 = _GEN_349 & ~_T_1463;
  assign stopEn134 = _GEN_349 & ~_T_1489;
  assign stopEn135 = _GEN_349 & ~_T_1396;
  assign stopEn136 = _GEN_349 & ~_T_1400;
  assign stopEn137 = _GEN_349 & ~_T_1403;
  assign stopEn138 = _GEN_349 & ~_T_1503;
  assign stopEn139 = _GEN_361 & ~_T_1393;
  assign stopEn140 = _GEN_361 & ~_T_1396;
  assign stopEn141 = _GEN_361 & ~_T_1403;
  assign stopEn142 = _GEN_361 & ~_T_1595;
  assign stopEn143 = _GEN_369 & ~_T_1393;
  assign stopEn144 = _GEN_369 & ~_T_1396;
  assign stopEn145 = _GEN_369 & ~_T_1403;
  assign stopEn146 = _GEN_369 & ~_T_1595;
  assign stopEn147 = _GEN_377 & ~_T_1393;
  assign stopEn148 = _GEN_377 & ~_T_1396;
  assign stopEn149 = _GEN_377 & ~_T_1403;
  assign stopEn150 = _GEN_377 & ~_T_1595;
  assign stopEn151 = _T_1663 & ~_T_1666;
  assign stopEn152 = _T_1663 & ~_T_1670;
  assign stopEn153 = _T_1663 & ~_T_1674;
  assign stopEn154 = _T_1663 & ~_T_1678;
  assign stopEn155 = _T_1663 & ~_T_1682;
  assign stopEn156 = _T_1712 & ~_T_1715;
  assign stopEn157 = _T_1712 & ~_T_1719;
  assign stopEn158 = _T_1712 & ~_T_1723;
  assign stopEn159 = _T_1712 & ~_T_1727;
  assign stopEn160 = _T_1712 & ~_T_1731;
  assign stopEn161 = _T_1712 & ~_T_1735;
  assign stopEn162 = _T_1765 & ~_T_1768;
  assign stopEn163 = _T_1765 & ~_T_1772;
  assign stopEn164 = _T_1765 & ~_T_1776;
  assign stopEn165 = _T_1765 & ~_T_1780;
  assign stopEn166 = _T_1765 & ~_T_1784;
  assign stopEn167 = _T_1813 & ~_T_1816;
  assign stopEn168 = _T_1813 & ~_T_1820;
  assign stopEn169 = _T_1813 & ~_T_1824;
  assign stopEn170 = _T_1813 & ~_T_1828;
  assign stopEn171 = _T_1813 & ~_T_1832;
  assign stopEn172 = _T_1892 & ~_T_1907;
  assign stopEn173 = _T_1931 & ~_T_1941;
  assign stopEn174 = _T_1931 & ~_T_1954;
  assign stopEn175 = _T_1931 & ~_T_1961;
  assign stopEn176 = _T_1969 & ~_T_1973;
  assign stopEn177 = ~_T_1980;
  assign stopEn178 = _T_2033 & ~_T_2039;
  assign stopEn179 = _T_2042 & ~_T_2050;
  assign TLMonitor_37_or63 = stopEn0 | stopEn1;
  assign TLMonitor_37_or130 = stopEn3 | stopEn4;
  assign TLMonitor_37_or64 = stopEn2 | TLMonitor_37_or130;
  assign TLMonitor_37_or31 = TLMonitor_37_or63 | TLMonitor_37_or64;
  assign TLMonitor_37_or132 = stopEn6 | stopEn7;
  assign TLMonitor_37_or65 = stopEn5 | TLMonitor_37_or132;
  assign TLMonitor_37_or134 = stopEn9 | stopEn10;
  assign TLMonitor_37_or66 = stopEn8 | TLMonitor_37_or134;
  assign TLMonitor_37_or32 = TLMonitor_37_or65 | TLMonitor_37_or66;
  assign TLMonitor_37_or15 = TLMonitor_37_or31 | TLMonitor_37_or32;
  assign TLMonitor_37_or67 = stopEn11 | stopEn12;
  assign TLMonitor_37_or138 = stopEn14 | stopEn15;
  assign TLMonitor_37_or68 = stopEn13 | TLMonitor_37_or138;
  assign TLMonitor_37_or33 = TLMonitor_37_or67 | TLMonitor_37_or68;
  assign TLMonitor_37_or140 = stopEn17 | stopEn18;
  assign TLMonitor_37_or69 = stopEn16 | TLMonitor_37_or140;
  assign TLMonitor_37_or142 = stopEn20 | stopEn21;
  assign TLMonitor_37_or70 = stopEn19 | TLMonitor_37_or142;
  assign TLMonitor_37_or34 = TLMonitor_37_or69 | TLMonitor_37_or70;
  assign TLMonitor_37_or16 = TLMonitor_37_or33 | TLMonitor_37_or34;
  assign TLMonitor_37_or7 = TLMonitor_37_or15 | TLMonitor_37_or16;
  assign TLMonitor_37_or71 = stopEn22 | stopEn23;
  assign TLMonitor_37_or146 = stopEn25 | stopEn26;
  assign TLMonitor_37_or72 = stopEn24 | TLMonitor_37_or146;
  assign TLMonitor_37_or35 = TLMonitor_37_or71 | TLMonitor_37_or72;
  assign TLMonitor_37_or148 = stopEn28 | stopEn29;
  assign TLMonitor_37_or73 = stopEn27 | TLMonitor_37_or148;
  assign TLMonitor_37_or150 = stopEn31 | stopEn32;
  assign TLMonitor_37_or74 = stopEn30 | TLMonitor_37_or150;
  assign TLMonitor_37_or36 = TLMonitor_37_or73 | TLMonitor_37_or74;
  assign TLMonitor_37_or17 = TLMonitor_37_or35 | TLMonitor_37_or36;
  assign TLMonitor_37_or152 = stopEn34 | stopEn35;
  assign TLMonitor_37_or75 = stopEn33 | TLMonitor_37_or152;
  assign TLMonitor_37_or154 = stopEn37 | stopEn38;
  assign TLMonitor_37_or76 = stopEn36 | TLMonitor_37_or154;
  assign TLMonitor_37_or37 = TLMonitor_37_or75 | TLMonitor_37_or76;
  assign TLMonitor_37_or156 = stopEn40 | stopEn41;
  assign TLMonitor_37_or77 = stopEn39 | TLMonitor_37_or156;
  assign TLMonitor_37_or158 = stopEn43 | stopEn44;
  assign TLMonitor_37_or78 = stopEn42 | TLMonitor_37_or158;
  assign TLMonitor_37_or38 = TLMonitor_37_or77 | TLMonitor_37_or78;
  assign TLMonitor_37_or18 = TLMonitor_37_or37 | TLMonitor_37_or38;
  assign TLMonitor_37_or8 = TLMonitor_37_or17 | TLMonitor_37_or18;
  assign TLMonitor_37_or3 = TLMonitor_37_or7 | TLMonitor_37_or8;
  assign TLMonitor_37_or79 = stopEn45 | stopEn46;
  assign TLMonitor_37_or162 = stopEn48 | stopEn49;
  assign TLMonitor_37_or80 = stopEn47 | TLMonitor_37_or162;
  assign TLMonitor_37_or39 = TLMonitor_37_or79 | TLMonitor_37_or80;
  assign TLMonitor_37_or164 = stopEn51 | stopEn52;
  assign TLMonitor_37_or81 = stopEn50 | TLMonitor_37_or164;
  assign TLMonitor_37_or166 = stopEn54 | stopEn55;
  assign TLMonitor_37_or82 = stopEn53 | TLMonitor_37_or166;
  assign TLMonitor_37_or40 = TLMonitor_37_or81 | TLMonitor_37_or82;
  assign TLMonitor_37_or19 = TLMonitor_37_or39 | TLMonitor_37_or40;
  assign TLMonitor_37_or83 = stopEn56 | stopEn57;
  assign TLMonitor_37_or170 = stopEn59 | stopEn60;
  assign TLMonitor_37_or84 = stopEn58 | TLMonitor_37_or170;
  assign TLMonitor_37_or41 = TLMonitor_37_or83 | TLMonitor_37_or84;
  assign TLMonitor_37_or172 = stopEn62 | stopEn63;
  assign TLMonitor_37_or85 = stopEn61 | TLMonitor_37_or172;
  assign TLMonitor_37_or174 = stopEn65 | stopEn66;
  assign TLMonitor_37_or86 = stopEn64 | TLMonitor_37_or174;
  assign TLMonitor_37_or42 = TLMonitor_37_or85 | TLMonitor_37_or86;
  assign TLMonitor_37_or20 = TLMonitor_37_or41 | TLMonitor_37_or42;
  assign TLMonitor_37_or9 = TLMonitor_37_or19 | TLMonitor_37_or20;
  assign TLMonitor_37_or87 = stopEn67 | stopEn68;
  assign TLMonitor_37_or178 = stopEn70 | stopEn71;
  assign TLMonitor_37_or88 = stopEn69 | TLMonitor_37_or178;
  assign TLMonitor_37_or43 = TLMonitor_37_or87 | TLMonitor_37_or88;
  assign TLMonitor_37_or180 = stopEn73 | stopEn74;
  assign TLMonitor_37_or89 = stopEn72 | TLMonitor_37_or180;
  assign TLMonitor_37_or182 = stopEn76 | stopEn77;
  assign TLMonitor_37_or90 = stopEn75 | TLMonitor_37_or182;
  assign TLMonitor_37_or44 = TLMonitor_37_or89 | TLMonitor_37_or90;
  assign TLMonitor_37_or21 = TLMonitor_37_or43 | TLMonitor_37_or44;
  assign TLMonitor_37_or184 = stopEn79 | stopEn80;
  assign TLMonitor_37_or91 = stopEn78 | TLMonitor_37_or184;
  assign TLMonitor_37_or186 = stopEn82 | stopEn83;
  assign TLMonitor_37_or92 = stopEn81 | TLMonitor_37_or186;
  assign TLMonitor_37_or45 = TLMonitor_37_or91 | TLMonitor_37_or92;
  assign TLMonitor_37_or188 = stopEn85 | stopEn86;
  assign TLMonitor_37_or93 = stopEn84 | TLMonitor_37_or188;
  assign TLMonitor_37_or190 = stopEn88 | stopEn89;
  assign TLMonitor_37_or94 = stopEn87 | TLMonitor_37_or190;
  assign TLMonitor_37_or46 = TLMonitor_37_or93 | TLMonitor_37_or94;
  assign TLMonitor_37_or22 = TLMonitor_37_or45 | TLMonitor_37_or46;
  assign TLMonitor_37_or10 = TLMonitor_37_or21 | TLMonitor_37_or22;
  assign TLMonitor_37_or4 = TLMonitor_37_or9 | TLMonitor_37_or10;
  assign TLMonitor_37_or1 = TLMonitor_37_or3 | TLMonitor_37_or4;
  assign TLMonitor_37_or95 = stopEn90 | stopEn91;
  assign TLMonitor_37_or194 = stopEn93 | stopEn94;
  assign TLMonitor_37_or96 = stopEn92 | TLMonitor_37_or194;
  assign TLMonitor_37_or47 = TLMonitor_37_or95 | TLMonitor_37_or96;
  assign TLMonitor_37_or196 = stopEn96 | stopEn97;
  assign TLMonitor_37_or97 = stopEn95 | TLMonitor_37_or196;
  assign TLMonitor_37_or198 = stopEn99 | stopEn100;
  assign TLMonitor_37_or98 = stopEn98 | TLMonitor_37_or198;
  assign TLMonitor_37_or48 = TLMonitor_37_or97 | TLMonitor_37_or98;
  assign TLMonitor_37_or23 = TLMonitor_37_or47 | TLMonitor_37_or48;
  assign TLMonitor_37_or99 = stopEn101 | stopEn102;
  assign TLMonitor_37_or202 = stopEn104 | stopEn105;
  assign TLMonitor_37_or100 = stopEn103 | TLMonitor_37_or202;
  assign TLMonitor_37_or49 = TLMonitor_37_or99 | TLMonitor_37_or100;
  assign TLMonitor_37_or204 = stopEn107 | stopEn108;
  assign TLMonitor_37_or101 = stopEn106 | TLMonitor_37_or204;
  assign TLMonitor_37_or206 = stopEn110 | stopEn111;
  assign TLMonitor_37_or102 = stopEn109 | TLMonitor_37_or206;
  assign TLMonitor_37_or50 = TLMonitor_37_or101 | TLMonitor_37_or102;
  assign TLMonitor_37_or24 = TLMonitor_37_or49 | TLMonitor_37_or50;
  assign TLMonitor_37_or11 = TLMonitor_37_or23 | TLMonitor_37_or24;
  assign TLMonitor_37_or103 = stopEn112 | stopEn113;
  assign TLMonitor_37_or210 = stopEn115 | stopEn116;
  assign TLMonitor_37_or104 = stopEn114 | TLMonitor_37_or210;
  assign TLMonitor_37_or51 = TLMonitor_37_or103 | TLMonitor_37_or104;
  assign TLMonitor_37_or212 = stopEn118 | stopEn119;
  assign TLMonitor_37_or105 = stopEn117 | TLMonitor_37_or212;
  assign TLMonitor_37_or214 = stopEn121 | stopEn122;
  assign TLMonitor_37_or106 = stopEn120 | TLMonitor_37_or214;
  assign TLMonitor_37_or52 = TLMonitor_37_or105 | TLMonitor_37_or106;
  assign TLMonitor_37_or25 = TLMonitor_37_or51 | TLMonitor_37_or52;
  assign TLMonitor_37_or216 = stopEn124 | stopEn125;
  assign TLMonitor_37_or107 = stopEn123 | TLMonitor_37_or216;
  assign TLMonitor_37_or218 = stopEn127 | stopEn128;
  assign TLMonitor_37_or108 = stopEn126 | TLMonitor_37_or218;
  assign TLMonitor_37_or53 = TLMonitor_37_or107 | TLMonitor_37_or108;
  assign TLMonitor_37_or220 = stopEn130 | stopEn131;
  assign TLMonitor_37_or109 = stopEn129 | TLMonitor_37_or220;
  assign TLMonitor_37_or222 = stopEn133 | stopEn134;
  assign TLMonitor_37_or110 = stopEn132 | TLMonitor_37_or222;
  assign TLMonitor_37_or54 = TLMonitor_37_or109 | TLMonitor_37_or110;
  assign TLMonitor_37_or26 = TLMonitor_37_or53 | TLMonitor_37_or54;
  assign TLMonitor_37_or12 = TLMonitor_37_or25 | TLMonitor_37_or26;
  assign TLMonitor_37_or5 = TLMonitor_37_or11 | TLMonitor_37_or12;
  assign TLMonitor_37_or111 = stopEn135 | stopEn136;
  assign TLMonitor_37_or226 = stopEn138 | stopEn139;
  assign TLMonitor_37_or112 = stopEn137 | TLMonitor_37_or226;
  assign TLMonitor_37_or55 = TLMonitor_37_or111 | TLMonitor_37_or112;
  assign TLMonitor_37_or228 = stopEn141 | stopEn142;
  assign TLMonitor_37_or113 = stopEn140 | TLMonitor_37_or228;
  assign TLMonitor_37_or230 = stopEn144 | stopEn145;
  assign TLMonitor_37_or114 = stopEn143 | TLMonitor_37_or230;
  assign TLMonitor_37_or56 = TLMonitor_37_or113 | TLMonitor_37_or114;
  assign TLMonitor_37_or27 = TLMonitor_37_or55 | TLMonitor_37_or56;
  assign TLMonitor_37_or115 = stopEn146 | stopEn147;
  assign TLMonitor_37_or234 = stopEn149 | stopEn150;
  assign TLMonitor_37_or116 = stopEn148 | TLMonitor_37_or234;
  assign TLMonitor_37_or57 = TLMonitor_37_or115 | TLMonitor_37_or116;
  assign TLMonitor_37_or236 = stopEn152 | stopEn153;
  assign TLMonitor_37_or117 = stopEn151 | TLMonitor_37_or236;
  assign TLMonitor_37_or238 = stopEn155 | stopEn156;
  assign TLMonitor_37_or118 = stopEn154 | TLMonitor_37_or238;
  assign TLMonitor_37_or58 = TLMonitor_37_or117 | TLMonitor_37_or118;
  assign TLMonitor_37_or28 = TLMonitor_37_or57 | TLMonitor_37_or58;
  assign TLMonitor_37_or13 = TLMonitor_37_or27 | TLMonitor_37_or28;
  assign TLMonitor_37_or119 = stopEn157 | stopEn158;
  assign TLMonitor_37_or242 = stopEn160 | stopEn161;
  assign TLMonitor_37_or120 = stopEn159 | TLMonitor_37_or242;
  assign TLMonitor_37_or59 = TLMonitor_37_or119 | TLMonitor_37_or120;
  assign TLMonitor_37_or244 = stopEn163 | stopEn164;
  assign TLMonitor_37_or121 = stopEn162 | TLMonitor_37_or244;
  assign TLMonitor_37_or246 = stopEn166 | stopEn167;
  assign TLMonitor_37_or122 = stopEn165 | TLMonitor_37_or246;
  assign TLMonitor_37_or60 = TLMonitor_37_or121 | TLMonitor_37_or122;
  assign TLMonitor_37_or29 = TLMonitor_37_or59 | TLMonitor_37_or60;
  assign TLMonitor_37_or248 = stopEn169 | stopEn170;
  assign TLMonitor_37_or123 = stopEn168 | TLMonitor_37_or248;
  assign TLMonitor_37_or250 = stopEn172 | stopEn173;
  assign TLMonitor_37_or124 = stopEn171 | TLMonitor_37_or250;
  assign TLMonitor_37_or61 = TLMonitor_37_or123 | TLMonitor_37_or124;
  assign TLMonitor_37_or252 = stopEn175 | stopEn176;
  assign TLMonitor_37_or125 = stopEn174 | TLMonitor_37_or252;
  assign TLMonitor_37_or254 = stopEn178 | stopEn179;
  assign TLMonitor_37_or126 = stopEn177 | TLMonitor_37_or254;
  assign TLMonitor_37_or62 = TLMonitor_37_or125 | TLMonitor_37_or126;
  assign TLMonitor_37_or30 = TLMonitor_37_or61 | TLMonitor_37_or62;
  assign TLMonitor_37_or14 = TLMonitor_37_or29 | TLMonitor_37_or30;
  assign TLMonitor_37_or6 = TLMonitor_37_or13 | TLMonitor_37_or14;
  assign TLMonitor_37_or2 = TLMonitor_37_or5 | TLMonitor_37_or6;
  assign TLMonitor_37_or0 = TLMonitor_37_or1 | TLMonitor_37_or2;
  assign metaAssert = TLMonitor_37_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1646 = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1657 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1658 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1659 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1660 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1661 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1694 = _RAND_6[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1705 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1706 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1707 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1708 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_1709 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1710 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_1748 = _RAND_13[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_1759 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_1760 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1761 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_1762 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_1763 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_1796 = _RAND_19[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_1807 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_1808 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_1809 = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_1810 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_1811 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  inflight = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  inflight_opcodes = _RAND_26[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  inflight_sizes = _RAND_27[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_1845 = _RAND_28[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_1863 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_2006 = _RAND_30[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_2015 = _RAND_31[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  TLMonitor_37_metaAssert = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_1646 <= 9'h0;
    end else if (reset) begin
      _T_1646 <= 9'h0;
    end else if (_T_1637) begin
      if (_T_1649) begin
        if (~io_in_a_bits_opcode[2]) begin
          _T_1646 <= _T_1642;
        end else begin
          _T_1646 <= 9'h0;
        end
      end else begin
        _T_1646 <= _T_1648;
      end
    end
    if (metaReset) begin
      _T_1657 <= 3'h0;
    end else if (_T_1685) begin
      _T_1657 <= io_in_a_bits_opcode;
    end
    if (metaReset) begin
      _T_1658 <= 3'h0;
    end else if (_T_1685) begin
      _T_1658 <= io_in_a_bits_param;
    end
    if (metaReset) begin
      _T_1659 <= 4'h0;
    end else if (_T_1685) begin
      _T_1659 <= io_in_a_bits_size;
    end
    if (metaReset) begin
      _T_1660 <= 2'h0;
    end else if (_T_1685) begin
      _T_1660 <= io_in_a_bits_source;
    end
    if (metaReset) begin
      _T_1661 <= 32'h0;
    end else if (_T_1685) begin
      _T_1661 <= io_in_a_bits_address;
    end
    if (metaReset) begin
      _T_1694 <= 9'h0;
    end else if (reset) begin
      _T_1694 <= 9'h0;
    end else if (_T_1686) begin
      if (_T_1697) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1694 <= _T_1691;
        end else begin
          _T_1694 <= 9'h0;
        end
      end else begin
        _T_1694 <= _T_1696;
      end
    end
    if (metaReset) begin
      _T_1705 <= 3'h0;
    end else if (_T_1738) begin
      _T_1705 <= io_in_d_bits_opcode;
    end
    if (metaReset) begin
      _T_1706 <= 2'h0;
    end else if (_T_1738) begin
      _T_1706 <= io_in_d_bits_param;
    end
    if (metaReset) begin
      _T_1707 <= 4'h0;
    end else if (_T_1738) begin
      _T_1707 <= io_in_d_bits_size;
    end
    if (metaReset) begin
      _T_1708 <= 2'h0;
    end else if (_T_1738) begin
      _T_1708 <= io_in_d_bits_source;
    end
    if (metaReset) begin
      _T_1709 <= 2'h0;
    end else if (_T_1738) begin
      _T_1709 <= io_in_d_bits_sink;
    end
    if (metaReset) begin
      _T_1710 <= 1'h0;
    end else if (_T_1738) begin
      _T_1710 <= io_in_d_bits_denied;
    end
    if (metaReset) begin
      _T_1748 <= 9'h0;
    end else if (reset) begin
      _T_1748 <= 9'h0;
    end else if (_T_1739) begin
      if (_T_1751) begin
        _T_1748 <= 9'h0;
      end else begin
        _T_1748 <= _T_1750;
      end
    end
    if (metaReset) begin
      _T_1759 <= 3'h0;
    end else if (_T_1787) begin
      _T_1759 <= io_in_b_bits_opcode;
    end
    if (metaReset) begin
      _T_1760 <= 2'h0;
    end else if (_T_1787) begin
      _T_1760 <= io_in_b_bits_param;
    end
    if (metaReset) begin
      _T_1761 <= 4'h0;
    end else if (_T_1787) begin
      _T_1761 <= io_in_b_bits_size;
    end
    if (metaReset) begin
      _T_1762 <= 2'h0;
    end else if (_T_1787) begin
      _T_1762 <= io_in_b_bits_source;
    end
    if (metaReset) begin
      _T_1763 <= 32'h0;
    end else if (_T_1787) begin
      _T_1763 <= io_in_b_bits_address;
    end
    if (metaReset) begin
      _T_1796 <= 9'h0;
    end else if (reset) begin
      _T_1796 <= 9'h0;
    end else if (_T_1788) begin
      if (_T_1799) begin
        if (io_in_c_bits_opcode[0]) begin
          _T_1796 <= _T_1793;
        end else begin
          _T_1796 <= 9'h0;
        end
      end else begin
        _T_1796 <= _T_1798;
      end
    end
    if (metaReset) begin
      _T_1807 <= 3'h0;
    end else if (_T_1835) begin
      _T_1807 <= io_in_c_bits_opcode;
    end
    if (metaReset) begin
      _T_1808 <= 3'h0;
    end else if (_T_1835) begin
      _T_1808 <= io_in_c_bits_param;
    end
    if (metaReset) begin
      _T_1809 <= 4'h0;
    end else if (_T_1835) begin
      _T_1809 <= io_in_c_bits_size;
    end
    if (metaReset) begin
      _T_1810 <= 2'h0;
    end else if (_T_1835) begin
      _T_1810 <= io_in_c_bits_source;
    end
    if (metaReset) begin
      _T_1811 <= 32'h0;
    end else if (_T_1835) begin
      _T_1811 <= io_in_c_bits_address;
    end
    if (metaReset) begin
      inflight <= 3'h0;
    end else if (reset) begin
      inflight <= 3'h0;
    end else begin
      inflight <= _T_1984;
    end
    if (metaReset) begin
      inflight_opcodes <= 12'h0;
    end else if (reset) begin
      inflight_opcodes <= 12'h0;
    end else begin
      inflight_opcodes <= _T_1987;
    end
    if (metaReset) begin
      inflight_sizes <= 24'h0;
    end else if (reset) begin
      inflight_sizes <= 24'h0;
    end else begin
      inflight_sizes <= _T_1990;
    end
    if (metaReset) begin
      _T_1845 <= 9'h0;
    end else if (reset) begin
      _T_1845 <= 9'h0;
    end else if (_T_1637) begin
      if (a_first) begin
        if (~io_in_a_bits_opcode[2]) begin
          _T_1845 <= _T_1642;
        end else begin
          _T_1845 <= 9'h0;
        end
      end else begin
        _T_1845 <= _T_1847;
      end
    end
    if (metaReset) begin
      _T_1863 <= 9'h0;
    end else if (reset) begin
      _T_1863 <= 9'h0;
    end else if (_T_1686) begin
      if (d_first) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1863 <= _T_1691;
        end else begin
          _T_1863 <= 9'h0;
        end
      end else begin
        _T_1863 <= _T_1865;
      end
    end
    if (metaReset) begin
      _T_2006 <= 4'h0;
    end else if (reset) begin
      _T_2006 <= 4'h0;
    end else begin
      _T_2006 <= _T_2054;
    end
    if (metaReset) begin
      _T_2015 <= 9'h0;
    end else if (reset) begin
      _T_2015 <= 9'h0;
    end else if (_T_1686) begin
      if (_T_2018) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_2015 <= _T_1691;
        end else begin
          _T_2015 <= 9'h0;
        end
      end else begin
        _T_2015 <= _T_2017;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & ~_T_141) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & ~_T_141) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & ~_T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & ~_T_167) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & ~_T_170) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & ~_T_170) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & ~_T_174) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & ~_T_174) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & ~_T_177) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & ~_T_177) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & ~_T_181) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & ~_T_181) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & ~_T_186) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & ~_T_186) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & ~_T_190) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & ~_T_190) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_141) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_141) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_167) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_170) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_170) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_174) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_174) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_177) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_177) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_181) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_181) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_268) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_268) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_186) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_186) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_190) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_190) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & ~_T_344) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type which is unexpected using diplomatic parameters\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & ~_T_344) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & ~_T_170) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & ~_T_170) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & ~_T_177) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & ~_T_177) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & ~_T_354) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & ~_T_354) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & ~_T_358) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & ~_T_358) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & ~_T_190) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & ~_T_190) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & ~_T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & ~_T_436) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & ~_T_170) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & ~_T_170) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & ~_T_177) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & ~_T_177) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & ~_T_354) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & ~_T_354) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & ~_T_358) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & ~_T_358) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & ~_T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & ~_T_436) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & ~_T_170) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & ~_T_170) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & ~_T_177) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & ~_T_177) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & ~_T_354) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & ~_T_354) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & ~_T_540) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & ~_T_540) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_592) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_592) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_170) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_170) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_177) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_177) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_602) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_602) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_358) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_358) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_592) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_592) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_170) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_170) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_177) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_177) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_668) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_668) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_358) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_358) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & ~_T_736) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & ~_T_736) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & ~_T_170) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID\nThe diplomacy information for the edge is as follows:\nMaster Name = Core 0 DCache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(0,1)\n\nMaster Name = Core 0 DCache MMIO\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(1,2)\n\nMaster Name = Core 0 ICache\nvisibility = List(AddressSet(0x0, ~0x0))\nemits = acquireT = TransferSizes[1, 4096]\nacquireB = TransferSizes[1, 4096]\narithmetic = TransferSizes[1, 4096]\nlogical = TransferSizes[1, 4096]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\nsourceId = IdRange(2,3)\n\n\nSlave Port Beatbytes = 8\nSlave Port MinLatency = 3\n\nSlave Name = error\nSlave Address = List(AddressSet(0x3000, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 4096]\nputFull = TransferSizes[1, 4096]\nputPartial = TransferSizes[1, 4096]\nhint = TransferSizes[1, 4096]\n\n\n\nSlave Name = plic\nSlave Address = List(AddressSet(0xc000000, 0x3ffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = clint\nSlave Address = List(AddressSet(0x2000000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = dmInner\nSlave Address = List(AddressSet(0x0, 0xfff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[1, 8]\nlogical = TransferSizes[1, 8]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = bootrom\nSlave Address = List(AddressSet(0x10000, 0xffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[0, 0]\nputPartial = TransferSizes[0, 0]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x80000000, 0xfffffff))\nsupports = acquireT = TransferSizes[1, 64]\nacquireB = TransferSizes[1, 64]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 64]\nputPartial = TransferSizes[1, 64]\nhint = TransferSizes[0, 0]\n\n\n\nSlave Name = ldut\nSlave Address = List(AddressSet(0x60000000, 0x1fffffff))\nsupports = acquireT = TransferSizes[0, 0]\nacquireB = TransferSizes[0, 0]\narithmetic = TransferSizes[0, 0]\nlogical = TransferSizes[0, 0]\nget = TransferSizes[1, 64]\nputFull = TransferSizes[1, 256]\nputPartial = TransferSizes[1, 256]\nhint = TransferSizes[0, 0]\n\n\n\n\n (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & ~_T_170) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & ~_T_177) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & ~_T_177) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & ~_T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid opcode param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & ~_T_746) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & ~_T_358) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & ~_T_358) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & ~_T_190) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & ~_T_190) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~_T_758) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~_T_758) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & ~_T_769) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & ~_T_769) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & ~_T_773) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & ~_T_773) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & ~_T_777) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & ~_T_777) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & ~_T_781) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & ~_T_781) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & ~_T_785) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & ~_T_785) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_769) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_769) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_773) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_773) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_800) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_800) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_804) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_804) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_781) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_781) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & ~_T_769) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & ~_T_769) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & ~_T_773) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & ~_T_773) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & ~_T_800) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & ~_T_800) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & ~_T_804) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & ~_T_804) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & ~_T_837) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & ~_T_837) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & ~_T_769) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & ~_T_769) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & ~_T_777) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & ~_T_777) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & ~_T_781) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & ~_T_781) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & ~_T_769) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & ~_T_769) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & ~_T_777) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & ~_T_777) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & ~_T_837) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & ~_T_837) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & ~_T_769) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & ~_T_769) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & ~_T_777) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & ~_T_777) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & ~_T_781) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & ~_T_781) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & ~_T_898) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & ~_T_898) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_1077) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type which is unexpected using diplomatic parameters (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_1077) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_1090) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_1090) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_1094) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_1098) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_1098) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type which is unexpected using diplomatic parameters (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & ~reset) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & ~_T_1127) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & ~_T_1127) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & ~_T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & ~_T_1094) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & ~_T_1098) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & ~_T_1098) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type which is unexpected using diplomatic parameters (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & ~reset) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & ~_T_1127) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & ~_T_1127) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & ~_T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & ~_T_1094) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & ~reset) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & ~_T_1127) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & ~_T_1127) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & ~_T_1203) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & ~_T_1203) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by master (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~reset) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1094) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & ~reset) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & ~_T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & ~_T_1094) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & ~reset) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & ~_T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & ~_T_1094) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & ~_T_1098) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & ~_T_1098) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1393) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1393) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1396) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1396) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1400) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1400) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1403) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1403) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1407) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1407) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & ~_T_1393) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & ~_T_1393) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & ~_T_1396) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & ~_T_1396) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & ~_T_1400) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & ~_T_1400) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & ~_T_1403) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & ~_T_1403) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & ~_T_1407) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & ~_T_1407) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & ~_T_1463) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & ~_T_1463) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & ~_T_1489) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & ~_T_1489) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & ~_T_1396) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & ~_T_1396) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & ~_T_1400) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & ~_T_1400) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & ~_T_1403) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & ~_T_1403) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & ~_T_1503) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & ~_T_1503) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & ~_T_1463) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & ~_T_1463) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & ~_T_1489) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & ~_T_1489) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & ~_T_1396) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & ~_T_1396) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & ~_T_1400) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & ~_T_1400) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & ~_T_1403) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & ~_T_1403) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & ~_T_1503) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & ~_T_1503) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & ~_T_1393) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & ~_T_1393) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & ~_T_1396) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & ~_T_1396) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & ~_T_1403) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & ~_T_1403) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & ~_T_1595) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & ~_T_1595) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_369 & ~_T_1393) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_369 & ~_T_1393) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_369 & ~_T_1396) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_369 & ~_T_1396) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_369 & ~_T_1403) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_369 & ~_T_1403) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_369 & ~_T_1595) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_369 & ~_T_1595) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_377 & ~_T_1393) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_377 & ~_T_1393) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_377 & ~_T_1396) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_377 & ~_T_1396) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_377 & ~_T_1403) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_377 & ~_T_1403) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_377 & ~_T_1595) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_377 & ~_T_1595) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1663 & ~_T_1666) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1663 & ~_T_1666) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1663 & ~_T_1670) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1663 & ~_T_1670) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1663 & ~_T_1674) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1663 & ~_T_1674) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1663 & ~_T_1678) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1663 & ~_T_1678) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1663 & ~_T_1682) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1663 & ~_T_1682) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1712 & ~_T_1715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1712 & ~_T_1715) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1712 & ~_T_1719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1712 & ~_T_1719) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1712 & ~_T_1723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1712 & ~_T_1723) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1712 & ~_T_1727) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1712 & ~_T_1727) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1712 & ~_T_1731) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1712 & ~_T_1731) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1712 & ~_T_1735) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1712 & ~_T_1735) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1765 & ~_T_1768) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1765 & ~_T_1768) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1765 & ~_T_1772) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1765 & ~_T_1772) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1765 & ~_T_1776) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1765 & ~_T_1776) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1765 & ~_T_1780) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1765 & ~_T_1780) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1765 & ~_T_1784) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1765 & ~_T_1784) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1813 & ~_T_1816) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1813 & ~_T_1816) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1813 & ~_T_1820) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1813 & ~_T_1820) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1813 & ~_T_1824) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1813 & ~_T_1824) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1813 & ~_T_1828) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1813 & ~_T_1828) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1813 & ~_T_1832) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1813 & ~_T_1832) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1892 & ~_T_1907) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1892 & ~_T_1907) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1931 & ~_T_1941) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1931 & ~_T_1941) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1931 & ~_T_1954) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1931 & ~_T_1954) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1931 & ~_T_1961) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1931 & ~_T_1961) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1969 & ~_T_1973) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1969 & ~_T_1973) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1980) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1980) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2033 & ~_T_2039) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2033 & ~_T_2039) begin
          $fatal; // @[Monitor.scala 51:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2042 & ~_T_2050) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2042 & ~_T_2050) begin
          $fatal; // @[Monitor.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    if (metaReset) begin
      TLMonitor_37_metaAssert <= 1'h0;
    end else begin
      TLMonitor_37_metaAssert <= TLMonitor_37_metaAssert | TLMonitor_37_or0;
    end
  end
endmodule
module Queue_32(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input  [63:0] io_enq_bits_data,
  input         io_enq_bits_corrupt,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_corrupt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_15_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_5_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_1;
  wire [2:0] ram_param__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_param__T_15_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_param__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_param__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_param__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_param__T_5_en; // @[Decoupled.scala 218:16]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_2;
  wire [3:0] ram_size__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_size__T_15_addr; // @[Decoupled.scala 218:16]
  wire [3:0] ram_size__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_size__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_size__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_size__T_5_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_source [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_3;
  wire [1:0] ram_source__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_source__T_15_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_source__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_source__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_source__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_source__T_5_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_address [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_4;
  wire [31:0] ram_address__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_address__T_15_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_address__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_address__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_address__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_address__T_5_en; // @[Decoupled.scala 218:16]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_5;
  wire [7:0] ram_mask__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_mask__T_15_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_mask__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_mask__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_mask__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_mask__T_5_en; // @[Decoupled.scala 218:16]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16]
  reg [63:0] _RAND_6;
  wire [63:0] ram_data__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_data__T_15_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_data__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_data__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_data__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_data__T_5_en; // @[Decoupled.scala 218:16]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_7;
  wire  ram_corrupt__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_15_addr; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_en; // @[Decoupled.scala 218:16]
  reg  _T; // @[Counter.scala 29:33]
  reg [31:0] _RAND_8;
  reg  _T_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_9;
  reg  maybe_full; // @[Decoupled.scala 221:27]
  reg [31:0] _RAND_10;
  wire  ptr_match; // @[Decoupled.scala 223:33]
  wire  empty; // @[Decoupled.scala 224:25]
  wire  full; // @[Decoupled.scala 225:24]
  wire  do_enq; // @[Decoupled.scala 40:37]
  wire  do_deq; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Counter.scala 39:22]
  wire  _T_11; // @[Counter.scala 39:22]
  wire  _T_12; // @[Decoupled.scala 236:16]
  wire [29:0] Queue_32_covSum;
  assign ram_opcode__T_15_addr = _T_1;
  assign ram_opcode__T_15_data = ram_opcode[ram_opcode__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_opcode__T_5_data = io_enq_bits_opcode;
  assign ram_opcode__T_5_addr = _T;
  assign ram_opcode__T_5_mask = 1'h1;
  assign ram_opcode__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_param__T_15_addr = _T_1;
  assign ram_param__T_15_data = ram_param[ram_param__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_param__T_5_data = io_enq_bits_param;
  assign ram_param__T_5_addr = _T;
  assign ram_param__T_5_mask = 1'h1;
  assign ram_param__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_size__T_15_addr = _T_1;
  assign ram_size__T_15_data = ram_size[ram_size__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_size__T_5_data = io_enq_bits_size;
  assign ram_size__T_5_addr = _T;
  assign ram_size__T_5_mask = 1'h1;
  assign ram_size__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_source__T_15_addr = _T_1;
  assign ram_source__T_15_data = ram_source[ram_source__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_source__T_5_data = io_enq_bits_source;
  assign ram_source__T_5_addr = _T;
  assign ram_source__T_5_mask = 1'h1;
  assign ram_source__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_address__T_15_addr = _T_1;
  assign ram_address__T_15_data = ram_address[ram_address__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_address__T_5_data = io_enq_bits_address;
  assign ram_address__T_5_addr = _T;
  assign ram_address__T_5_mask = 1'h1;
  assign ram_address__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_mask__T_15_addr = _T_1;
  assign ram_mask__T_15_data = ram_mask[ram_mask__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_mask__T_5_data = io_enq_bits_mask;
  assign ram_mask__T_5_addr = _T;
  assign ram_mask__T_5_mask = 1'h1;
  assign ram_mask__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_15_addr = _T_1;
  assign ram_data__T_15_data = ram_data[ram_data__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_data__T_5_data = io_enq_bits_data;
  assign ram_data__T_5_addr = _T;
  assign ram_data__T_5_mask = 1'h1;
  assign ram_data__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt__T_15_addr = _T_1;
  assign ram_corrupt__T_15_data = ram_corrupt[ram_corrupt__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_corrupt__T_5_data = io_enq_bits_corrupt;
  assign ram_corrupt__T_5_addr = _T;
  assign ram_corrupt__T_5_mask = 1'h1;
  assign ram_corrupt__T_5_en = io_enq_ready & io_enq_valid;
  assign ptr_match = _T == _T_1; // @[Decoupled.scala 223:33]
  assign empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  assign full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  assign do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = _T + 1'h1; // @[Counter.scala 39:22]
  assign _T_11 = _T_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_12 = do_enq != do_deq; // @[Decoupled.scala 236:16]
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:16]
  assign io_deq_bits_opcode = ram_opcode__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_param = ram_param__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_size = ram_size__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_source = ram_source__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_address = ram_address__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_mask = ram_mask__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_data = ram_data__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_corrupt = ram_corrupt__T_15_data; // @[Decoupled.scala 242:15]
  assign Queue_32_covSum = 30'h0;
  assign io_covSum = Queue_32_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_opcode__T_5_en & ram_opcode__T_5_mask) begin
      ram_opcode[ram_opcode__T_5_addr] <= ram_opcode__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_param__T_5_en & ram_param__T_5_mask) begin
      ram_param[ram_param__T_5_addr] <= ram_param__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_size__T_5_en & ram_size__T_5_mask) begin
      ram_size[ram_size__T_5_addr] <= ram_size__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_source__T_5_en & ram_source__T_5_mask) begin
      ram_source[ram_source__T_5_addr] <= ram_source__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_address__T_5_en & ram_address__T_5_mask) begin
      ram_address[ram_address__T_5_addr] <= ram_address__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_mask__T_5_en & ram_mask__T_5_mask) begin
      ram_mask[ram_mask__T_5_addr] <= ram_mask__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_data__T_5_en & ram_data__T_5_mask) begin
      ram_data[ram_data__T_5_addr] <= ram_data__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_corrupt__T_5_en & ram_corrupt__T_5_mask) begin
      ram_corrupt[ram_corrupt__T_5_addr] <= ram_corrupt__T_5_data; // @[Decoupled.scala 218:16]
    end
    if (metaReset) begin
      _T <= 1'h0;
    end else if (reset) begin
      _T <= 1'h0;
    end else if (do_enq) begin
      _T <= _T_8;
    end
    if (metaReset) begin
      _T_1 <= 1'h0;
    end else if (reset) begin
      _T_1 <= 1'h0;
    end else if (do_deq) begin
      _T_1 <= _T_11;
    end
    if (metaReset) begin
      maybe_full <= 1'h0;
    end else if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_12) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_33(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_source,
  input  [1:0]  io_enq_bits_sink,
  input         io_enq_bits_denied,
  input  [63:0] io_enq_bits_data,
  input         io_enq_bits_corrupt,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_source,
  output [1:0]  io_deq_bits_sink,
  output        io_deq_bits_denied,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_corrupt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_15_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_5_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_param [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_1;
  wire [1:0] ram_param__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_param__T_15_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_param__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_param__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_param__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_param__T_5_en; // @[Decoupled.scala 218:16]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_2;
  wire [3:0] ram_size__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_size__T_15_addr; // @[Decoupled.scala 218:16]
  wire [3:0] ram_size__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_size__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_size__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_size__T_5_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_source [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_3;
  wire [1:0] ram_source__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_source__T_15_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_source__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_source__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_source__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_source__T_5_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_sink [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_4;
  wire [1:0] ram_sink__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_sink__T_15_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_sink__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_sink__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_sink__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_sink__T_5_en; // @[Decoupled.scala 218:16]
  reg  ram_denied [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_5;
  wire  ram_denied__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_denied__T_15_addr; // @[Decoupled.scala 218:16]
  wire  ram_denied__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_denied__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_denied__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_denied__T_5_en; // @[Decoupled.scala 218:16]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16]
  reg [63:0] _RAND_6;
  wire [63:0] ram_data__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_data__T_15_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_data__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_data__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_data__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_data__T_5_en; // @[Decoupled.scala 218:16]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_7;
  wire  ram_corrupt__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_15_addr; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_en; // @[Decoupled.scala 218:16]
  reg  _T; // @[Counter.scala 29:33]
  reg [31:0] _RAND_8;
  reg  _T_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_9;
  reg  maybe_full; // @[Decoupled.scala 221:27]
  reg [31:0] _RAND_10;
  wire  ptr_match; // @[Decoupled.scala 223:33]
  wire  empty; // @[Decoupled.scala 224:25]
  wire  full; // @[Decoupled.scala 225:24]
  wire  do_enq; // @[Decoupled.scala 40:37]
  wire  do_deq; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Counter.scala 39:22]
  wire  _T_11; // @[Counter.scala 39:22]
  wire  _T_12; // @[Decoupled.scala 236:16]
  wire [29:0] Queue_33_covSum;
  assign ram_opcode__T_15_addr = _T_1;
  assign ram_opcode__T_15_data = ram_opcode[ram_opcode__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_opcode__T_5_data = io_enq_bits_opcode;
  assign ram_opcode__T_5_addr = _T;
  assign ram_opcode__T_5_mask = 1'h1;
  assign ram_opcode__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_param__T_15_addr = _T_1;
  assign ram_param__T_15_data = ram_param[ram_param__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_param__T_5_data = io_enq_bits_param;
  assign ram_param__T_5_addr = _T;
  assign ram_param__T_5_mask = 1'h1;
  assign ram_param__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_size__T_15_addr = _T_1;
  assign ram_size__T_15_data = ram_size[ram_size__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_size__T_5_data = io_enq_bits_size;
  assign ram_size__T_5_addr = _T;
  assign ram_size__T_5_mask = 1'h1;
  assign ram_size__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_source__T_15_addr = _T_1;
  assign ram_source__T_15_data = ram_source[ram_source__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_source__T_5_data = io_enq_bits_source;
  assign ram_source__T_5_addr = _T;
  assign ram_source__T_5_mask = 1'h1;
  assign ram_source__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_sink__T_15_addr = _T_1;
  assign ram_sink__T_15_data = ram_sink[ram_sink__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_sink__T_5_data = io_enq_bits_sink;
  assign ram_sink__T_5_addr = _T;
  assign ram_sink__T_5_mask = 1'h1;
  assign ram_sink__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_denied__T_15_addr = _T_1;
  assign ram_denied__T_15_data = ram_denied[ram_denied__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_denied__T_5_data = io_enq_bits_denied;
  assign ram_denied__T_5_addr = _T;
  assign ram_denied__T_5_mask = 1'h1;
  assign ram_denied__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_15_addr = _T_1;
  assign ram_data__T_15_data = ram_data[ram_data__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_data__T_5_data = io_enq_bits_data;
  assign ram_data__T_5_addr = _T;
  assign ram_data__T_5_mask = 1'h1;
  assign ram_data__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt__T_15_addr = _T_1;
  assign ram_corrupt__T_15_data = ram_corrupt[ram_corrupt__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_corrupt__T_5_data = io_enq_bits_corrupt;
  assign ram_corrupt__T_5_addr = _T;
  assign ram_corrupt__T_5_mask = 1'h1;
  assign ram_corrupt__T_5_en = io_enq_ready & io_enq_valid;
  assign ptr_match = _T == _T_1; // @[Decoupled.scala 223:33]
  assign empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  assign full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  assign do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = _T + 1'h1; // @[Counter.scala 39:22]
  assign _T_11 = _T_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_12 = do_enq != do_deq; // @[Decoupled.scala 236:16]
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:16]
  assign io_deq_bits_opcode = ram_opcode__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_param = ram_param__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_size = ram_size__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_source = ram_source__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_sink = ram_sink__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_denied = ram_denied__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_data = ram_data__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_corrupt = ram_corrupt__T_15_data; // @[Decoupled.scala 242:15]
  assign Queue_33_covSum = 30'h0;
  assign io_covSum = Queue_33_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_opcode__T_5_en & ram_opcode__T_5_mask) begin
      ram_opcode[ram_opcode__T_5_addr] <= ram_opcode__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_param__T_5_en & ram_param__T_5_mask) begin
      ram_param[ram_param__T_5_addr] <= ram_param__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_size__T_5_en & ram_size__T_5_mask) begin
      ram_size[ram_size__T_5_addr] <= ram_size__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_source__T_5_en & ram_source__T_5_mask) begin
      ram_source[ram_source__T_5_addr] <= ram_source__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_sink__T_5_en & ram_sink__T_5_mask) begin
      ram_sink[ram_sink__T_5_addr] <= ram_sink__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_denied__T_5_en & ram_denied__T_5_mask) begin
      ram_denied[ram_denied__T_5_addr] <= ram_denied__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_data__T_5_en & ram_data__T_5_mask) begin
      ram_data[ram_data__T_5_addr] <= ram_data__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_corrupt__T_5_en & ram_corrupt__T_5_mask) begin
      ram_corrupt[ram_corrupt__T_5_addr] <= ram_corrupt__T_5_data; // @[Decoupled.scala 218:16]
    end
    if (metaReset) begin
      _T <= 1'h0;
    end else if (reset) begin
      _T <= 1'h0;
    end else if (do_enq) begin
      _T <= _T_8;
    end
    if (metaReset) begin
      _T_1 <= 1'h0;
    end else if (reset) begin
      _T_1 <= 1'h0;
    end else if (do_deq) begin
      _T_1 <= _T_11;
    end
    if (metaReset) begin
      maybe_full <= 1'h0;
    end else if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_12) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_34(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input         io_enq_bits_corrupt,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output        io_deq_bits_corrupt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_15_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_5_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_param [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_1;
  wire [1:0] ram_param__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_param__T_15_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_param__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_param__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_param__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_param__T_5_en; // @[Decoupled.scala 218:16]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_2;
  wire [3:0] ram_size__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_size__T_15_addr; // @[Decoupled.scala 218:16]
  wire [3:0] ram_size__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_size__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_size__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_size__T_5_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_source [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_3;
  wire [1:0] ram_source__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_source__T_15_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_source__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_source__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_source__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_source__T_5_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_address [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_4;
  wire [31:0] ram_address__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_address__T_15_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_address__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_address__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_address__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_address__T_5_en; // @[Decoupled.scala 218:16]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_5;
  wire [7:0] ram_mask__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_mask__T_15_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_mask__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_mask__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_mask__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_mask__T_5_en; // @[Decoupled.scala 218:16]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_6;
  wire  ram_corrupt__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_15_addr; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_en; // @[Decoupled.scala 218:16]
  reg  _T; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  reg  _T_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_8;
  reg  maybe_full; // @[Decoupled.scala 221:27]
  reg [31:0] _RAND_9;
  wire  ptr_match; // @[Decoupled.scala 223:33]
  wire  empty; // @[Decoupled.scala 224:25]
  wire  full; // @[Decoupled.scala 225:24]
  wire  do_enq; // @[Decoupled.scala 40:37]
  wire  do_deq; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Counter.scala 39:22]
  wire  _T_11; // @[Counter.scala 39:22]
  wire  _T_12; // @[Decoupled.scala 236:16]
  wire [29:0] Queue_34_covSum;
  assign ram_opcode__T_15_addr = _T_1;
  assign ram_opcode__T_15_data = ram_opcode[ram_opcode__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_opcode__T_5_data = io_enq_bits_opcode;
  assign ram_opcode__T_5_addr = _T;
  assign ram_opcode__T_5_mask = 1'h1;
  assign ram_opcode__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_param__T_15_addr = _T_1;
  assign ram_param__T_15_data = ram_param[ram_param__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_param__T_5_data = io_enq_bits_param;
  assign ram_param__T_5_addr = _T;
  assign ram_param__T_5_mask = 1'h1;
  assign ram_param__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_size__T_15_addr = _T_1;
  assign ram_size__T_15_data = ram_size[ram_size__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_size__T_5_data = io_enq_bits_size;
  assign ram_size__T_5_addr = _T;
  assign ram_size__T_5_mask = 1'h1;
  assign ram_size__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_source__T_15_addr = _T_1;
  assign ram_source__T_15_data = ram_source[ram_source__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_source__T_5_data = io_enq_bits_source;
  assign ram_source__T_5_addr = _T;
  assign ram_source__T_5_mask = 1'h1;
  assign ram_source__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_address__T_15_addr = _T_1;
  assign ram_address__T_15_data = ram_address[ram_address__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_address__T_5_data = io_enq_bits_address;
  assign ram_address__T_5_addr = _T;
  assign ram_address__T_5_mask = 1'h1;
  assign ram_address__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_mask__T_15_addr = _T_1;
  assign ram_mask__T_15_data = ram_mask[ram_mask__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_mask__T_5_data = io_enq_bits_mask;
  assign ram_mask__T_5_addr = _T;
  assign ram_mask__T_5_mask = 1'h1;
  assign ram_mask__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt__T_15_addr = _T_1;
  assign ram_corrupt__T_15_data = ram_corrupt[ram_corrupt__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_corrupt__T_5_data = io_enq_bits_corrupt;
  assign ram_corrupt__T_5_addr = _T;
  assign ram_corrupt__T_5_mask = 1'h1;
  assign ram_corrupt__T_5_en = io_enq_ready & io_enq_valid;
  assign ptr_match = _T == _T_1; // @[Decoupled.scala 223:33]
  assign empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  assign full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  assign do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = _T + 1'h1; // @[Counter.scala 39:22]
  assign _T_11 = _T_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_12 = do_enq != do_deq; // @[Decoupled.scala 236:16]
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:16]
  assign io_deq_bits_opcode = ram_opcode__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_param = ram_param__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_size = ram_size__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_source = ram_source__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_address = ram_address__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_mask = ram_mask__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_corrupt = ram_corrupt__T_15_data; // @[Decoupled.scala 242:15]
  assign Queue_34_covSum = 30'h0;
  assign io_covSum = Queue_34_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_6[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  maybe_full = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_opcode__T_5_en & ram_opcode__T_5_mask) begin
      ram_opcode[ram_opcode__T_5_addr] <= ram_opcode__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_param__T_5_en & ram_param__T_5_mask) begin
      ram_param[ram_param__T_5_addr] <= ram_param__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_size__T_5_en & ram_size__T_5_mask) begin
      ram_size[ram_size__T_5_addr] <= ram_size__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_source__T_5_en & ram_source__T_5_mask) begin
      ram_source[ram_source__T_5_addr] <= ram_source__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_address__T_5_en & ram_address__T_5_mask) begin
      ram_address[ram_address__T_5_addr] <= ram_address__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_mask__T_5_en & ram_mask__T_5_mask) begin
      ram_mask[ram_mask__T_5_addr] <= ram_mask__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_corrupt__T_5_en & ram_corrupt__T_5_mask) begin
      ram_corrupt[ram_corrupt__T_5_addr] <= ram_corrupt__T_5_data; // @[Decoupled.scala 218:16]
    end
    if (metaReset) begin
      _T <= 1'h0;
    end else if (reset) begin
      _T <= 1'h0;
    end else if (do_enq) begin
      _T <= _T_8;
    end
    if (metaReset) begin
      _T_1 <= 1'h0;
    end else if (reset) begin
      _T_1 <= 1'h0;
    end else if (do_deq) begin
      _T_1 <= _T_11;
    end
    if (metaReset) begin
      maybe_full <= 1'h0;
    end else if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_12) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_35(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_corrupt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_15_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_opcode__T_5_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_1;
  wire [2:0] ram_param__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_param__T_15_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_param__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_param__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_param__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_param__T_5_en; // @[Decoupled.scala 218:16]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_2;
  wire [3:0] ram_size__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_size__T_15_addr; // @[Decoupled.scala 218:16]
  wire [3:0] ram_size__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_size__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_size__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_size__T_5_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_source [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_3;
  wire [1:0] ram_source__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_source__T_15_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_source__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_source__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_source__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_source__T_5_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_address [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_4;
  wire [31:0] ram_address__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_address__T_15_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_address__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_address__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_address__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_address__T_5_en; // @[Decoupled.scala 218:16]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16]
  reg [63:0] _RAND_5;
  wire [63:0] ram_data__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_data__T_15_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_data__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_data__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_data__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_data__T_5_en; // @[Decoupled.scala 218:16]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_6;
  wire  ram_corrupt__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_15_addr; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_corrupt__T_5_en; // @[Decoupled.scala 218:16]
  reg  _T; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  reg  _T_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_8;
  reg  maybe_full; // @[Decoupled.scala 221:27]
  reg [31:0] _RAND_9;
  wire  ptr_match; // @[Decoupled.scala 223:33]
  wire  empty; // @[Decoupled.scala 224:25]
  wire  full; // @[Decoupled.scala 225:24]
  wire  do_enq; // @[Decoupled.scala 40:37]
  wire  do_deq; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Counter.scala 39:22]
  wire  _T_11; // @[Counter.scala 39:22]
  wire  _T_12; // @[Decoupled.scala 236:16]
  wire [29:0] Queue_35_covSum;
  assign ram_opcode__T_15_addr = _T_1;
  assign ram_opcode__T_15_data = ram_opcode[ram_opcode__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_opcode__T_5_data = io_enq_bits_opcode;
  assign ram_opcode__T_5_addr = _T;
  assign ram_opcode__T_5_mask = 1'h1;
  assign ram_opcode__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_param__T_15_addr = _T_1;
  assign ram_param__T_15_data = ram_param[ram_param__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_param__T_5_data = io_enq_bits_param;
  assign ram_param__T_5_addr = _T;
  assign ram_param__T_5_mask = 1'h1;
  assign ram_param__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_size__T_15_addr = _T_1;
  assign ram_size__T_15_data = ram_size[ram_size__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_size__T_5_data = io_enq_bits_size;
  assign ram_size__T_5_addr = _T;
  assign ram_size__T_5_mask = 1'h1;
  assign ram_size__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_source__T_15_addr = _T_1;
  assign ram_source__T_15_data = ram_source[ram_source__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_source__T_5_data = io_enq_bits_source;
  assign ram_source__T_5_addr = _T;
  assign ram_source__T_5_mask = 1'h1;
  assign ram_source__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_address__T_15_addr = _T_1;
  assign ram_address__T_15_data = ram_address[ram_address__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_address__T_5_data = io_enq_bits_address;
  assign ram_address__T_5_addr = _T;
  assign ram_address__T_5_mask = 1'h1;
  assign ram_address__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_15_addr = _T_1;
  assign ram_data__T_15_data = ram_data[ram_data__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_data__T_5_data = io_enq_bits_data;
  assign ram_data__T_5_addr = _T;
  assign ram_data__T_5_mask = 1'h1;
  assign ram_data__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt__T_15_addr = _T_1;
  assign ram_corrupt__T_15_data = ram_corrupt[ram_corrupt__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_corrupt__T_5_data = 1'h0;
  assign ram_corrupt__T_5_addr = _T;
  assign ram_corrupt__T_5_mask = 1'h1;
  assign ram_corrupt__T_5_en = io_enq_ready & io_enq_valid;
  assign ptr_match = _T == _T_1; // @[Decoupled.scala 223:33]
  assign empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  assign full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  assign do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = _T + 1'h1; // @[Counter.scala 39:22]
  assign _T_11 = _T_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_12 = do_enq != do_deq; // @[Decoupled.scala 236:16]
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:16]
  assign io_deq_bits_opcode = ram_opcode__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_param = ram_param__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_size = ram_size__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_source = ram_source__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_address = ram_address__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_data = ram_data__T_15_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_corrupt = ram_corrupt__T_15_data; // @[Decoupled.scala 242:15]
  assign Queue_35_covSum = 30'h0;
  assign io_covSum = Queue_35_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_5[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_6[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  maybe_full = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_opcode__T_5_en & ram_opcode__T_5_mask) begin
      ram_opcode[ram_opcode__T_5_addr] <= ram_opcode__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_param__T_5_en & ram_param__T_5_mask) begin
      ram_param[ram_param__T_5_addr] <= ram_param__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_size__T_5_en & ram_size__T_5_mask) begin
      ram_size[ram_size__T_5_addr] <= ram_size__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_source__T_5_en & ram_source__T_5_mask) begin
      ram_source[ram_source__T_5_addr] <= ram_source__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_address__T_5_en & ram_address__T_5_mask) begin
      ram_address[ram_address__T_5_addr] <= ram_address__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_data__T_5_en & ram_data__T_5_mask) begin
      ram_data[ram_data__T_5_addr] <= ram_data__T_5_data; // @[Decoupled.scala 218:16]
    end
    if(ram_corrupt__T_5_en & ram_corrupt__T_5_mask) begin
      ram_corrupt[ram_corrupt__T_5_addr] <= ram_corrupt__T_5_data; // @[Decoupled.scala 218:16]
    end
    if (metaReset) begin
      _T <= 1'h0;
    end else if (reset) begin
      _T <= 1'h0;
    end else if (do_enq) begin
      _T <= _T_8;
    end
    if (metaReset) begin
      _T_1 <= 1'h0;
    end else if (reset) begin
      _T_1 <= 1'h0;
    end else if (do_deq) begin
      _T_1 <= _T_11;
    end
    if (metaReset) begin
      maybe_full <= 1'h0;
    end else if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_12) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_36(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_sink,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [1:0] ram_sink [0:1]; // @[Decoupled.scala 218:16]
  reg [31:0] _RAND_0;
  wire [1:0] ram_sink__T_15_data; // @[Decoupled.scala 218:16]
  wire  ram_sink__T_15_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_sink__T_5_data; // @[Decoupled.scala 218:16]
  wire  ram_sink__T_5_addr; // @[Decoupled.scala 218:16]
  wire  ram_sink__T_5_mask; // @[Decoupled.scala 218:16]
  wire  ram_sink__T_5_en; // @[Decoupled.scala 218:16]
  reg  _T; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg  _T_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  maybe_full; // @[Decoupled.scala 221:27]
  reg [31:0] _RAND_3;
  wire  ptr_match; // @[Decoupled.scala 223:33]
  wire  empty; // @[Decoupled.scala 224:25]
  wire  full; // @[Decoupled.scala 225:24]
  wire  do_enq; // @[Decoupled.scala 40:37]
  wire  do_deq; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Counter.scala 39:22]
  wire  _T_11; // @[Counter.scala 39:22]
  wire  _T_12; // @[Decoupled.scala 236:16]
  wire [29:0] Queue_36_covSum;
  assign ram_sink__T_15_addr = _T_1;
  assign ram_sink__T_15_data = ram_sink[ram_sink__T_15_addr]; // @[Decoupled.scala 218:16]
  assign ram_sink__T_5_data = io_enq_bits_sink;
  assign ram_sink__T_5_addr = _T;
  assign ram_sink__T_5_mask = 1'h1;
  assign ram_sink__T_5_en = io_enq_ready & io_enq_valid;
  assign ptr_match = _T == _T_1; // @[Decoupled.scala 223:33]
  assign empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  assign full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  assign do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = _T + 1'h1; // @[Counter.scala 39:22]
  assign _T_11 = _T_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_12 = do_enq != do_deq; // @[Decoupled.scala 236:16]
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:16]
  assign io_deq_bits_sink = ram_sink__T_15_data; // @[Decoupled.scala 242:15]
  assign Queue_36_covSum = 30'h0;
  assign io_covSum = Queue_36_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_sink__T_5_en & ram_sink__T_5_mask) begin
      ram_sink[ram_sink__T_5_addr] <= ram_sink__T_5_data; // @[Decoupled.scala 218:16]
    end
    if (metaReset) begin
      _T <= 1'h0;
    end else if (reset) begin
      _T <= 1'h0;
    end else if (do_enq) begin
      _T <= _T_8;
    end
    if (metaReset) begin
      _T_1 <= 1'h0;
    end else if (reset) begin
      _T_1 <= 1'h0;
    end else if (do_deq) begin
      _T_1 <= _T_11;
    end
    if (metaReset) begin
      maybe_full <= 1'h0;
    end else if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_12) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module SynchronizerShiftReg_w1_d3(
  input         clock,
  input         io_d,
  output        io_q,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         NonSyncResetSynchronizerPrimitiveShiftReg_d3_halt
);
  wire  NonSyncResetSynchronizerPrimitiveShiftReg_d3_clock; // @[ShiftReg.scala 45:23]
  wire  NonSyncResetSynchronizerPrimitiveShiftReg_d3_io_d; // @[ShiftReg.scala 45:23]
  wire  NonSyncResetSynchronizerPrimitiveShiftReg_d3_io_q; // @[ShiftReg.scala 45:23]
  wire [29:0] NonSyncResetSynchronizerPrimitiveShiftReg_d3_io_covSum; // @[ShiftReg.scala 45:23]
  wire  NonSyncResetSynchronizerPrimitiveShiftReg_d3_metaAssert; // @[ShiftReg.scala 45:23]
  wire  NonSyncResetSynchronizerPrimitiveShiftReg_d3_metaReset; // @[ShiftReg.scala 45:23]
  wire [29:0] SynchronizerShiftReg_w1_d3_covSum;
  wire [29:0] NonSyncResetSynchronizerPrimitiveShiftReg_d3_sum;
  wire  NonSyncResetSynchronizerPrimitiveShiftReg_d3_metaAssert_wire;
  NonSyncResetSynchronizerPrimitiveShiftReg_d3 NonSyncResetSynchronizerPrimitiveShiftReg_d3 ( // @[ShiftReg.scala 45:23]
    .clock(NonSyncResetSynchronizerPrimitiveShiftReg_d3_clock),
    .io_d(NonSyncResetSynchronizerPrimitiveShiftReg_d3_io_d),
    .io_q(NonSyncResetSynchronizerPrimitiveShiftReg_d3_io_q),
    .io_covSum(NonSyncResetSynchronizerPrimitiveShiftReg_d3_io_covSum),
    .metaAssert(NonSyncResetSynchronizerPrimitiveShiftReg_d3_metaAssert),
    .metaReset(NonSyncResetSynchronizerPrimitiveShiftReg_d3_metaReset)
  );
  assign io_q = NonSyncResetSynchronizerPrimitiveShiftReg_d3_io_q; // @[SynchronizerReg.scala 165:8]
  assign NonSyncResetSynchronizerPrimitiveShiftReg_d3_clock = clock;
  assign NonSyncResetSynchronizerPrimitiveShiftReg_d3_io_d = io_d; // @[ShiftReg.scala 47:16]
  assign SynchronizerShiftReg_w1_d3_covSum = 30'h0;
  assign NonSyncResetSynchronizerPrimitiveShiftReg_d3_sum = SynchronizerShiftReg_w1_d3_covSum + NonSyncResetSynchronizerPrimitiveShiftReg_d3_io_covSum;
  assign io_covSum = NonSyncResetSynchronizerPrimitiveShiftReg_d3_sum;
  assign NonSyncResetSynchronizerPrimitiveShiftReg_d3_metaAssert_wire = NonSyncResetSynchronizerPrimitiveShiftReg_d3_metaAssert;
  assign metaAssert = NonSyncResetSynchronizerPrimitiveShiftReg_d3_metaAssert_wire;
  assign NonSyncResetSynchronizerPrimitiveShiftReg_d3_metaReset = metaReset | NonSyncResetSynchronizerPrimitiveShiftReg_d3_halt;
endmodule
module FPUDecoder(
  input  [31:0] io_inst,
  output        io_sigs_wen,
  output        io_sigs_ren1,
  output        io_sigs_ren2,
  output        io_sigs_ren3,
  output        io_sigs_swap12,
  output        io_sigs_swap23,
  output        io_sigs_singleIn,
  output        io_sigs_singleOut,
  output        io_sigs_fromint,
  output        io_sigs_toint,
  output        io_sigs_fastpipe,
  output        io_sigs_fma,
  output        io_sigs_div,
  output        io_sigs_sqrt,
  output        io_sigs_wflags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [31:0] _T; // @[Decode.scala 14:65]
  wire [31:0] _T_2; // @[Decode.scala 14:65]
  wire  _T_3; // @[Decode.scala 14:121]
  wire [31:0] _T_4; // @[Decode.scala 14:65]
  wire  _T_5; // @[Decode.scala 14:121]
  wire [31:0] _T_6; // @[Decode.scala 14:65]
  wire  _T_7; // @[Decode.scala 14:121]
  wire  _T_9; // @[Decode.scala 15:30]
  wire [31:0] _T_10; // @[Decode.scala 14:65]
  wire  _T_11; // @[Decode.scala 14:121]
  wire [31:0] _T_12; // @[Decode.scala 14:65]
  wire  _T_13; // @[Decode.scala 14:121]
  wire [31:0] _T_14; // @[Decode.scala 14:65]
  wire  decoder_4; // @[Decode.scala 14:121]
  wire  _T_17; // @[Decode.scala 15:30]
  wire [31:0] _T_18; // @[Decode.scala 14:65]
  wire  _T_19; // @[Decode.scala 14:121]
  wire [31:0] _T_20; // @[Decode.scala 14:65]
  wire  _T_21; // @[Decode.scala 14:121]
  wire  _T_23; // @[Decode.scala 15:30]
  wire [31:0] _T_24; // @[Decode.scala 14:65]
  wire [31:0] _T_26; // @[Decode.scala 14:65]
  wire  _T_27; // @[Decode.scala 14:121]
  wire [31:0] _T_28; // @[Decode.scala 14:65]
  wire  _T_29; // @[Decode.scala 14:121]
  wire [31:0] _T_30; // @[Decode.scala 14:65]
  wire  _T_31; // @[Decode.scala 14:121]
  wire [31:0] _T_32; // @[Decode.scala 14:65]
  wire  _T_33; // @[Decode.scala 14:121]
  wire [31:0] _T_34; // @[Decode.scala 14:65]
  wire  _T_35; // @[Decode.scala 14:121]
  wire [31:0] _T_36; // @[Decode.scala 14:65]
  wire  _T_37; // @[Decode.scala 14:121]
  wire [31:0] _T_38; // @[Decode.scala 14:65]
  wire  _T_39; // @[Decode.scala 14:121]
  wire  _T_41; // @[Decode.scala 15:30]
  wire  _T_42; // @[Decode.scala 15:30]
  wire  _T_43; // @[Decode.scala 15:30]
  wire  _T_44; // @[Decode.scala 15:30]
  wire  _T_45; // @[Decode.scala 15:30]
  wire [31:0] _T_46; // @[Decode.scala 14:65]
  wire  _T_47; // @[Decode.scala 14:121]
  wire [31:0] _T_48; // @[Decode.scala 14:65]
  wire  _T_49; // @[Decode.scala 14:121]
  wire  _T_51; // @[Decode.scala 14:121]
  wire [31:0] _T_52; // @[Decode.scala 14:65]
  wire  _T_53; // @[Decode.scala 14:121]
  wire [31:0] _T_54; // @[Decode.scala 14:65]
  wire  _T_55; // @[Decode.scala 14:121]
  wire  _T_57; // @[Decode.scala 15:30]
  wire  _T_58; // @[Decode.scala 15:30]
  wire  _T_59; // @[Decode.scala 15:30]
  wire [31:0] _T_60; // @[Decode.scala 14:65]
  wire  _T_63; // @[Decode.scala 14:121]
  wire [31:0] _T_65; // @[Decode.scala 14:65]
  wire  _T_66; // @[Decode.scala 14:121]
  wire [31:0] _T_67; // @[Decode.scala 14:65]
  wire  _T_68; // @[Decode.scala 14:121]
  wire [31:0] _T_70; // @[Decode.scala 14:65]
  wire  _T_71; // @[Decode.scala 14:121]
  wire [31:0] _T_72; // @[Decode.scala 14:65]
  wire  _T_73; // @[Decode.scala 14:121]
  wire  _T_75; // @[Decode.scala 15:30]
  wire [31:0] _T_76; // @[Decode.scala 14:65]
  wire [31:0] _T_80; // @[Decode.scala 14:65]
  wire  _T_81; // @[Decode.scala 14:121]
  wire [31:0] _T_82; // @[Decode.scala 14:65]
  wire  _T_83; // @[Decode.scala 14:121]
  wire [31:0] _T_84; // @[Decode.scala 14:65]
  wire  _T_85; // @[Decode.scala 14:121]
  wire  _T_87; // @[Decode.scala 15:30]
  wire  _T_88; // @[Decode.scala 15:30]
  wire [29:0] FPUDecoder_covSum;
  assign _T = io_inst & 32'h40; // @[Decode.scala 14:65]
  assign _T_2 = io_inst & 32'h80000020; // @[Decode.scala 14:65]
  assign _T_3 = _T_2 == 32'h0; // @[Decode.scala 14:121]
  assign _T_4 = io_inst & 32'h30; // @[Decode.scala 14:65]
  assign _T_5 = _T_4 == 32'h0; // @[Decode.scala 14:121]
  assign _T_6 = io_inst & 32'h10000020; // @[Decode.scala 14:65]
  assign _T_7 = _T_6 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_9 = _T_3 | _T_5; // @[Decode.scala 15:30]
  assign _T_10 = io_inst & 32'h80000004; // @[Decode.scala 14:65]
  assign _T_11 = _T_10 == 32'h0; // @[Decode.scala 14:121]
  assign _T_12 = io_inst & 32'h10000004; // @[Decode.scala 14:65]
  assign _T_13 = _T_12 == 32'h0; // @[Decode.scala 14:121]
  assign _T_14 = io_inst & 32'h50; // @[Decode.scala 14:65]
  assign decoder_4 = _T_14 == 32'h40; // @[Decode.scala 14:121]
  assign _T_17 = _T_11 | _T_13; // @[Decode.scala 15:30]
  assign _T_18 = io_inst & 32'h40000004; // @[Decode.scala 14:65]
  assign _T_19 = _T_18 == 32'h0; // @[Decode.scala 14:121]
  assign _T_20 = io_inst & 32'h20; // @[Decode.scala 14:65]
  assign _T_21 = _T_20 == 32'h20; // @[Decode.scala 14:121]
  assign _T_23 = _T_19 | _T_21; // @[Decode.scala 15:30]
  assign _T_24 = io_inst & 32'h30000010; // @[Decode.scala 14:65]
  assign _T_26 = io_inst & 32'h82100020; // @[Decode.scala 14:65]
  assign _T_27 = _T_26 == 32'h0; // @[Decode.scala 14:121]
  assign _T_28 = io_inst & 32'h42000020; // @[Decode.scala 14:65]
  assign _T_29 = _T_28 == 32'h0; // @[Decode.scala 14:121]
  assign _T_30 = io_inst & 32'h2000030; // @[Decode.scala 14:65]
  assign _T_31 = _T_30 == 32'h0; // @[Decode.scala 14:121]
  assign _T_32 = io_inst & 32'h2103000; // @[Decode.scala 14:65]
  assign _T_33 = _T_32 == 32'h1000; // @[Decode.scala 14:121]
  assign _T_34 = io_inst & 32'h12002000; // @[Decode.scala 14:65]
  assign _T_35 = _T_34 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_36 = io_inst & 32'hd0100010; // @[Decode.scala 14:65]
  assign _T_37 = _T_36 == 32'h40000010; // @[Decode.scala 14:121]
  assign _T_38 = io_inst & 32'ha2000020; // @[Decode.scala 14:65]
  assign _T_39 = _T_38 == 32'h80000000; // @[Decode.scala 14:121]
  assign _T_41 = _T_27 | _T_29; // @[Decode.scala 15:30]
  assign _T_42 = _T_41 | _T_31; // @[Decode.scala 15:30]
  assign _T_43 = _T_42 | _T_33; // @[Decode.scala 15:30]
  assign _T_44 = _T_43 | _T_35; // @[Decode.scala 15:30]
  assign _T_45 = _T_44 | _T_37; // @[Decode.scala 15:30]
  assign _T_46 = io_inst & 32'h42001000; // @[Decode.scala 14:65]
  assign _T_47 = _T_46 == 32'h0; // @[Decode.scala 14:121]
  assign _T_48 = io_inst & 32'h22000004; // @[Decode.scala 14:65]
  assign _T_49 = _T_48 == 32'h0; // @[Decode.scala 14:121]
  assign _T_51 = _T_34 == 32'h0; // @[Decode.scala 14:121]
  assign _T_52 = io_inst & 32'h1040; // @[Decode.scala 14:65]
  assign _T_53 = _T_52 == 32'h0; // @[Decode.scala 14:121]
  assign _T_54 = io_inst & 32'h2000050; // @[Decode.scala 14:65]
  assign _T_55 = _T_54 == 32'h40; // @[Decode.scala 14:121]
  assign _T_57 = _T_47 | _T_49; // @[Decode.scala 15:30]
  assign _T_58 = _T_57 | _T_51; // @[Decode.scala 15:30]
  assign _T_59 = _T_58 | _T_53; // @[Decode.scala 15:30]
  assign _T_60 = io_inst & 32'h90000010; // @[Decode.scala 14:65]
  assign _T_63 = _T_60 == 32'h80000010; // @[Decode.scala 14:121]
  assign _T_65 = io_inst & 32'ha0000010; // @[Decode.scala 14:65]
  assign _T_66 = _T_65 == 32'h20000010; // @[Decode.scala 14:121]
  assign _T_67 = io_inst & 32'hd0000010; // @[Decode.scala 14:65]
  assign _T_68 = _T_67 == 32'h40000010; // @[Decode.scala 14:121]
  assign _T_70 = io_inst & 32'h70000004; // @[Decode.scala 14:65]
  assign _T_71 = _T_70 == 32'h0; // @[Decode.scala 14:121]
  assign _T_72 = io_inst & 32'h68000004; // @[Decode.scala 14:65]
  assign _T_73 = _T_72 == 32'h0; // @[Decode.scala 14:121]
  assign _T_75 = _T_71 | _T_73; // @[Decode.scala 15:30]
  assign _T_76 = io_inst & 32'h58000010; // @[Decode.scala 14:65]
  assign _T_80 = io_inst & 32'h20000004; // @[Decode.scala 14:65]
  assign _T_81 = _T_80 == 32'h0; // @[Decode.scala 14:121]
  assign _T_82 = io_inst & 32'h8002000; // @[Decode.scala 14:65]
  assign _T_83 = _T_82 == 32'h8000000; // @[Decode.scala 14:121]
  assign _T_84 = io_inst & 32'hc0000004; // @[Decode.scala 14:65]
  assign _T_85 = _T_84 == 32'h80000000; // @[Decode.scala 14:121]
  assign _T_87 = _T_81 | decoder_4; // @[Decode.scala 15:30]
  assign _T_88 = _T_87 | _T_83; // @[Decode.scala 15:30]
  assign io_sigs_wen = _T_9 | _T_7; // @[FPU.scala 135:40]
  assign io_sigs_ren1 = _T_17 | decoder_4; // @[FPU.scala 135:40]
  assign io_sigs_ren2 = _T_23 | decoder_4; // @[FPU.scala 135:40]
  assign io_sigs_ren3 = _T_14 == 32'h40; // @[FPU.scala 135:40]
  assign io_sigs_swap12 = _T == 32'h0; // @[FPU.scala 135:40]
  assign io_sigs_swap23 = _T_24 == 32'h10; // @[FPU.scala 135:40]
  assign io_sigs_singleIn = _T_45 | _T_39; // @[FPU.scala 135:40]
  assign io_sigs_singleOut = _T_59 | _T_55; // @[FPU.scala 135:40]
  assign io_sigs_fromint = _T_60 == 32'h90000010; // @[FPU.scala 135:40]
  assign io_sigs_toint = _T_21 | _T_63; // @[FPU.scala 135:40]
  assign io_sigs_fastpipe = _T_66 | _T_68; // @[FPU.scala 135:40]
  assign io_sigs_fma = _T_75 | decoder_4; // @[FPU.scala 135:40]
  assign io_sigs_div = _T_76 == 32'h18000010; // @[FPU.scala 135:40]
  assign io_sigs_sqrt = _T_67 == 32'h50000010; // @[FPU.scala 135:40]
  assign io_sigs_wflags = _T_88 | _T_85; // @[FPU.scala 135:40]
  assign FPUDecoder_covSum = 30'h0;
  assign io_covSum = FPUDecoder_covSum;
  assign metaAssert = 1'h0;
endmodule
module FPUFMAPipe(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_ren3,
  input         io_in_bits_swap23,
  input  [2:0]  io_in_bits_rm,
  input  [1:0]  io_in_bits_fmaCmd,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output [64:0] io_out_bits_data,
  output [4:0]  io_out_bits_exc,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         fma_halt
);
  wire  fma_clock; // @[FPU.scala 664:19]
  wire  fma_reset; // @[FPU.scala 664:19]
  wire  fma_io_validin; // @[FPU.scala 664:19]
  wire [1:0] fma_io_op; // @[FPU.scala 664:19]
  wire [32:0] fma_io_a; // @[FPU.scala 664:19]
  wire [32:0] fma_io_b; // @[FPU.scala 664:19]
  wire [32:0] fma_io_c; // @[FPU.scala 664:19]
  wire [2:0] fma_io_roundingMode; // @[FPU.scala 664:19]
  wire [32:0] fma_io_out; // @[FPU.scala 664:19]
  wire [4:0] fma_io_exceptionFlags; // @[FPU.scala 664:19]
  wire [29:0] fma_io_covSum; // @[FPU.scala 664:19]
  wire  fma_metaAssert; // @[FPU.scala 664:19]
  wire  fma_metaReset; // @[FPU.scala 664:19]
  reg  valid; // @[FPU.scala 652:18]
  reg [31:0] _RAND_0;
  reg [2:0] in_rm; // @[FPU.scala 653:15]
  reg [31:0] _RAND_1;
  reg [1:0] in_fmaCmd; // @[FPU.scala 653:15]
  reg [31:0] _RAND_2;
  reg [64:0] in_in1; // @[FPU.scala 653:15]
  reg [95:0] _RAND_3;
  reg [64:0] in_in2; // @[FPU.scala 653:15]
  reg [95:0] _RAND_4;
  reg [64:0] in_in3; // @[FPU.scala 653:15]
  reg [95:0] _RAND_5;
  wire [64:0] _T_1; // @[FPU.scala 656:32]
  wire [64:0] _T_3; // @[FPU.scala 656:50]
  wire  _T_4; // @[FPU.scala 661:21]
  wire [29:0] FPUFMAPipe_covSum;
  wire [29:0] fma_sum;
  wire  fma_metaAssert_wire;
  reg  FPUFMAPipe_metaAssert;
  reg [31:0] _RAND_6;
  MulAddRecFNPipe fma ( // @[FPU.scala 664:19]
    .clock(fma_clock),
    .reset(fma_reset),
    .io_validin(fma_io_validin),
    .io_op(fma_io_op),
    .io_a(fma_io_a),
    .io_b(fma_io_b),
    .io_c(fma_io_c),
    .io_roundingMode(fma_io_roundingMode),
    .io_out(fma_io_out),
    .io_exceptionFlags(fma_io_exceptionFlags),
    .io_covSum(fma_io_covSum),
    .metaAssert(fma_metaAssert),
    .metaReset(fma_metaReset)
  );
  assign _T_1 = io_in_bits_in1 ^ io_in_bits_in2; // @[FPU.scala 656:32]
  assign _T_3 = _T_1 & 65'h100000000; // @[FPU.scala 656:50]
  assign _T_4 = io_in_bits_ren3 | io_in_bits_swap23; // @[FPU.scala 661:21]
  assign io_out_bits_data = {{32'd0}, fma_io_out}; // @[FPU.scala 677:10]
  assign io_out_bits_exc = fma_io_exceptionFlags; // @[FPU.scala 677:10]
  assign fma_clock = clock;
  assign fma_reset = reset;
  assign fma_io_validin = valid; // @[FPU.scala 665:18]
  assign fma_io_op = in_fmaCmd; // @[FPU.scala 666:13]
  assign fma_io_a = in_in1[32:0]; // @[FPU.scala 669:12]
  assign fma_io_b = in_in2[32:0]; // @[FPU.scala 670:12]
  assign fma_io_c = in_in3[32:0]; // @[FPU.scala 671:12]
  assign fma_io_roundingMode = in_rm; // @[FPU.scala 667:23]
  assign FPUFMAPipe_covSum = 30'h0;
  assign fma_sum = FPUFMAPipe_covSum + fma_io_covSum;
  assign io_covSum = fma_sum;
  assign fma_metaAssert_wire = fma_metaAssert;
  assign metaAssert = FPUFMAPipe_metaAssert;
  assign fma_metaReset = metaReset | fma_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_rm = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_fmaCmd = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {3{`RANDOM}};
  in_in1 = _RAND_3[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {3{`RANDOM}};
  in_in2 = _RAND_4[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  in_in3 = _RAND_5[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  FPUFMAPipe_metaAssert = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      valid <= 1'h0;
    end else begin
      valid <= io_in_valid;
    end
    if (metaReset) begin
      in_rm <= 3'h0;
    end else if (io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      in_fmaCmd <= 2'h0;
    end else if (io_in_valid) begin
      in_fmaCmd <= io_in_bits_fmaCmd;
    end
    if (metaReset) begin
      in_in1 <= 65'h0;
    end else if (io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      in_in2 <= 65'h0;
    end else if (io_in_valid) begin
      if (io_in_bits_swap23) begin
        in_in2 <= 65'h80000000;
      end else begin
        in_in2 <= io_in_bits_in2;
      end
    end
    if (metaReset) begin
      in_in3 <= 65'h0;
    end else if (io_in_valid) begin
      if (~_T_4) begin
        in_in3 <= _T_3;
      end else begin
        in_in3 <= io_in_bits_in3;
      end
    end
    if (metaReset) begin
      FPUFMAPipe_metaAssert <= 1'h0;
    end else begin
      FPUFMAPipe_metaAssert <= FPUFMAPipe_metaAssert | fma_metaAssert_wire;
    end
  end
endmodule
module FPToInt(
  input         clock,
  input         io_in_valid,
  input         io_in_bits_ren2,
  input         io_in_bits_singleIn,
  input         io_in_bits_singleOut,
  input         io_in_bits_wflags,
  input  [2:0]  io_in_bits_rm,
  input  [1:0]  io_in_bits_typ,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  output [2:0]  io_out_bits_in_rm,
  output [64:0] io_out_bits_in_in1,
  output [64:0] io_out_bits_in_in2,
  output        io_out_bits_lt,
  output [63:0] io_out_bits_store,
  output [63:0] io_out_bits_toint,
  output [4:0]  io_out_bits_exc,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [64:0] dcmp_io_a; // @[FPU.scala 418:20]
  wire [64:0] dcmp_io_b; // @[FPU.scala 418:20]
  wire  dcmp_io_signaling; // @[FPU.scala 418:20]
  wire  dcmp_io_lt; // @[FPU.scala 418:20]
  wire  dcmp_io_eq; // @[FPU.scala 418:20]
  wire [4:0] dcmp_io_exceptionFlags; // @[FPU.scala 418:20]
  wire [29:0] dcmp_io_covSum; // @[FPU.scala 418:20]
  wire  dcmp_metaAssert; // @[FPU.scala 418:20]
  wire [64:0] RecFNToIN_io_in; // @[FPU.scala 445:24]
  wire [2:0] RecFNToIN_io_roundingMode; // @[FPU.scala 445:24]
  wire  RecFNToIN_io_signedOut; // @[FPU.scala 445:24]
  wire [63:0] RecFNToIN_io_out; // @[FPU.scala 445:24]
  wire [2:0] RecFNToIN_io_intExceptionFlags; // @[FPU.scala 445:24]
  wire [29:0] RecFNToIN_io_covSum; // @[FPU.scala 445:24]
  wire  RecFNToIN_metaAssert; // @[FPU.scala 445:24]
  wire [64:0] RecFNToIN_1_io_in; // @[FPU.scala 455:30]
  wire [2:0] RecFNToIN_1_io_roundingMode; // @[FPU.scala 455:30]
  wire  RecFNToIN_1_io_signedOut; // @[FPU.scala 455:30]
  wire [2:0] RecFNToIN_1_io_intExceptionFlags; // @[FPU.scala 455:30]
  wire [29:0] RecFNToIN_1_io_covSum; // @[FPU.scala 455:30]
  wire  RecFNToIN_1_metaAssert; // @[FPU.scala 455:30]
  reg  in_ren2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg  in_singleOut; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  in_wflags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [2:0] in_rm; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [1:0] in_typ; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [64:0] in_in1; // @[Reg.scala 15:16]
  reg [95:0] _RAND_5;
  reg [64:0] in_in2; // @[Reg.scala 15:16]
  reg [95:0] _RAND_6;
  wire  tag; // @[FPU.scala 423:13]
  wire  _T_4; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_6; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_9; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_12; // @[rawFloatFromRecFN.scala 56:33]
  wire [12:0] _T_14; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] _T_18; // @[Cat.scala 29:58]
  wire  _T_19; // @[fNFromRecFN.scala 50:39]
  wire [5:0] _T_22; // @[fNFromRecFN.scala 51:39]
  wire [52:0] _T_24; // @[fNFromRecFN.scala 52:42]
  wire [10:0] _T_28; // @[fNFromRecFN.scala 57:45]
  wire [10:0] _T_29; // @[fNFromRecFN.scala 55:16]
  wire  _T_30; // @[fNFromRecFN.scala 59:44]
  wire [10:0] _T_32; // @[Bitwise.scala 72:12]
  wire [10:0] _T_33; // @[fNFromRecFN.scala 59:15]
  wire [51:0] _T_35; // @[fNFromRecFN.scala 63:20]
  wire [51:0] _T_36; // @[fNFromRecFN.scala 61:16]
  wire [63:0] _T_38; // @[Cat.scala 29:58]
  wire [32:0] _T_43; // @[Cat.scala 29:58]
  wire  _T_46; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_48; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_51; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_54; // @[rawFloatFromRecFN.scala 56:33]
  wire [9:0] _T_56; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] _T_60; // @[Cat.scala 29:58]
  wire  _T_61; // @[fNFromRecFN.scala 50:39]
  wire [4:0] _T_64; // @[fNFromRecFN.scala 51:39]
  wire [23:0] _T_66; // @[fNFromRecFN.scala 52:42]
  wire [7:0] _T_70; // @[fNFromRecFN.scala 57:45]
  wire [7:0] _T_71; // @[fNFromRecFN.scala 55:16]
  wire  _T_72; // @[fNFromRecFN.scala 59:44]
  wire [7:0] _T_74; // @[Bitwise.scala 72:12]
  wire [7:0] _T_75; // @[fNFromRecFN.scala 59:15]
  wire [22:0] _T_77; // @[fNFromRecFN.scala 63:20]
  wire [22:0] _T_78; // @[fNFromRecFN.scala 61:16]
  wire [31:0] _T_80; // @[Cat.scala 29:58]
  wire  _T_83; // @[FPU.scala 203:56]
  wire [31:0] _T_85; // @[FPU.scala 394:44]
  wire [63:0] store; // @[Cat.scala 29:58]
  wire [63:0] _T_87; // @[Cat.scala 29:58]
  wire  _T_247; // @[FPU.scala 462:54]
  wire  _T_239; // @[FPU.scala 460:59]
  wire  _T_240; // @[FPU.scala 461:46]
  wire [30:0] _T_243; // @[Bitwise.scala 72:12]
  wire [63:0] _T_249; // @[Cat.scala 29:58]
  wire [63:0] _GEN_24; // @[FPU.scala 463:26]
  wire [63:0] _GEN_25; // @[FPU.scala 454:30]
  wire [1:0] _T_217; // @[Cat.scala 29:58]
  wire [2:0] _GEN_33; // @[FPU.scala 438:22]
  wire [2:0] _T_218; // @[FPU.scala 438:22]
  wire  _T_219; // @[FPU.scala 438:53]
  wire [63:0] _T_221; // @[FPU.scala 438:77]
  wire [63:0] _GEN_34; // @[FPU.scala 438:57]
  wire [63:0] _T_222; // @[FPU.scala 438:57]
  wire [63:0] _GEN_28; // @[FPU.scala 442:21]
  wire  _T_189; // @[FPU.scala 219:24]
  wire  _T_187; // @[FPU.scala 218:24]
  wire  _T_168; // @[FPU.scala 210:28]
  wire  _T_183; // @[FPU.scala 216:27]
  wire  _T_191; // @[FPU.scala 221:31]
  wire  _T_175; // @[FPU.scala 214:27]
  wire  _T_170; // @[FPU.scala 212:55]
  wire  _T_177; // @[FPU.scala 214:39]
  wire  _T_178; // @[FPU.scala 214:71]
  wire  _T_179; // @[FPU.scala 214:61]
  wire  _T_193; // @[FPU.scala 221:50]
  wire  _T_171; // @[FPU.scala 213:28]
  wire  _T_173; // @[FPU.scala 213:62]
  wire  _T_174; // @[FPU.scala 213:40]
  wire  _T_195; // @[FPU.scala 222:21]
  wire  _T_180; // @[FPU.scala 215:23]
  wire  _T_197; // @[FPU.scala 222:38]
  wire  _T_198; // @[FPU.scala 222:55]
  wire  _T_199; // @[FPU.scala 223:21]
  wire  _T_200; // @[FPU.scala 223:39]
  wire  _T_201; // @[FPU.scala 223:54]
  wire [9:0] _T_210; // @[Cat.scala 29:58]
  wire  _T_111; // @[FPU.scala 235:36]
  wire  _T_112; // @[FPU.scala 235:25]
  wire [11:0] _T_107; // @[FPU.scala 234:31]
  wire [11:0] _T_109; // @[FPU.scala 234:48]
  wire [8:0] _T_114; // @[Cat.scala 29:58]
  wire [8:0] _T_116; // @[FPU.scala 235:10]
  wire [75:0] _T_103; // @[FPU.scala 231:28]
  wire [32:0] _T_118; // @[Cat.scala 29:58]
  wire  _T_138; // @[FPU.scala 217:22]
  wire  _T_143; // @[FPU.scala 219:24]
  wire  _T_141; // @[FPU.scala 218:24]
  wire  _T_122; // @[FPU.scala 210:28]
  wire  _T_137; // @[FPU.scala 216:27]
  wire  _T_145; // @[FPU.scala 221:31]
  wire  _T_129; // @[FPU.scala 214:27]
  wire  _T_124; // @[FPU.scala 212:55]
  wire  _T_131; // @[FPU.scala 214:39]
  wire  _T_132; // @[FPU.scala 214:71]
  wire  _T_133; // @[FPU.scala 214:61]
  wire  _T_147; // @[FPU.scala 221:50]
  wire  _T_125; // @[FPU.scala 213:28]
  wire  _T_127; // @[FPU.scala 213:62]
  wire  _T_128; // @[FPU.scala 213:40]
  wire  _T_149; // @[FPU.scala 222:21]
  wire  _T_134; // @[FPU.scala 215:23]
  wire  _T_151; // @[FPU.scala 222:38]
  wire  _T_152; // @[FPU.scala 222:55]
  wire  _T_153; // @[FPU.scala 223:21]
  wire  _T_154; // @[FPU.scala 223:39]
  wire  _T_155; // @[FPU.scala 223:54]
  wire [9:0] _T_164; // @[Cat.scala 29:58]
  wire [9:0] _T_212; // @[package.scala 32:76]
  wire [63:0] _GEN_35; // @[FPU.scala 433:27]
  wire [63:0] _T_215; // @[FPU.scala 433:27]
  wire [63:0] _GEN_22; // @[FPU.scala 431:19]
  wire [63:0] toint; // @[FPU.scala 437:20]
  wire [31:0] _T_94; // @[Bitwise.scala 72:12]
  wire [63:0] _T_95; // @[Cat.scala 29:58]
  wire  _GEN_27; // @[FPU.scala 442:21]
  wire  _GEN_23; // @[FPU.scala 431:19]
  wire  intType; // @[FPU.scala 437:20]
  wire  _T_228; // @[FPU.scala 450:62]
  wire [4:0] _T_231; // @[Cat.scala 29:58]
  wire  _T_252; // @[FPU.scala 464:64]
  wire [4:0] _T_254; // @[Cat.scala 29:58]
  wire [4:0] _GEN_26; // @[FPU.scala 454:30]
  wire [4:0] _GEN_29; // @[FPU.scala 442:21]
  wire  _T_256; // @[FPU.scala 471:53]
  wire  _T_258; // @[FPU.scala 471:79]
  wire  _T_259; // @[FPU.scala 471:59]
  reg [4:0] FPToInt_state; // @[Register tracking FPToInt state]
  reg [31:0] _RAND_7;
  reg  FPToInt_cov [0:31]; // @[Coverage map for FPToInt]
  reg [31:0] _RAND_8;
  wire  FPToInt_cov_read_data; // @[Coverage map for FPToInt]
  wire [4:0] FPToInt_cov_read_addr; // @[Coverage map for FPToInt]
  wire  FPToInt_cov_write_data; // @[Coverage map for FPToInt]
  wire [4:0] FPToInt_cov_write_addr; // @[Coverage map for FPToInt]
  wire  FPToInt_cov_write_mask; // @[Coverage map for FPToInt]
  wire  FPToInt_cov_write_en; // @[Coverage map for FPToInt]
  reg [29:0] FPToInt_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_9;
  wire  in_wflags_shl;
  wire [4:0] in_wflags_pad;
  wire [1:0] in_singleOut_shl;
  wire [4:0] in_singleOut_pad;
  wire [3:0] in_typ_shl;
  wire [4:0] in_typ_pad;
  wire [4:0] in_ren2_shl;
  wire [4:0] in_ren2_pad;
  wire [4:0] FPToInt_xor1;
  wire [4:0] FPToInt_xor2;
  wire [4:0] FPToInt_xor0;
  wire [29:0] dcmp_sum;
  wire [29:0] RecFNToIN_sum;
  wire [29:0] RecFNToIN_1_sum;
  wire  dcmp_metaAssert_wire;
  wire  RecFNToIN_metaAssert_wire;
  wire  RecFNToIN_1_metaAssert_wire;
  wire  FPToInt_or2;
  wire  FPToInt_or0;
  CompareRecFN dcmp ( // @[FPU.scala 418:20]
    .io_a(dcmp_io_a),
    .io_b(dcmp_io_b),
    .io_signaling(dcmp_io_signaling),
    .io_lt(dcmp_io_lt),
    .io_eq(dcmp_io_eq),
    .io_exceptionFlags(dcmp_io_exceptionFlags),
    .io_covSum(dcmp_io_covSum),
    .metaAssert(dcmp_metaAssert)
  );
  RecFNToIN RecFNToIN ( // @[FPU.scala 445:24]
    .io_in(RecFNToIN_io_in),
    .io_roundingMode(RecFNToIN_io_roundingMode),
    .io_signedOut(RecFNToIN_io_signedOut),
    .io_out(RecFNToIN_io_out),
    .io_intExceptionFlags(RecFNToIN_io_intExceptionFlags),
    .io_covSum(RecFNToIN_io_covSum),
    .metaAssert(RecFNToIN_metaAssert)
  );
  RecFNToIN_1 RecFNToIN_1 ( // @[FPU.scala 455:30]
    .io_in(RecFNToIN_1_io_in),
    .io_roundingMode(RecFNToIN_1_io_roundingMode),
    .io_signedOut(RecFNToIN_1_io_signedOut),
    .io_intExceptionFlags(RecFNToIN_1_io_intExceptionFlags),
    .io_covSum(RecFNToIN_1_io_covSum),
    .metaAssert(RecFNToIN_1_metaAssert)
  );
  assign tag = ~in_singleOut; // @[FPU.scala 423:13]
  assign _T_4 = in_in1[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_6 = in_in1[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign _T_9 = _T_6 & in_in1[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign _T_12 = _T_6 & ~in_in1[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign _T_14 = {1'b0,$signed(in_in1[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign _T_18 = {1'h0,~_T_4,in_in1[51:0]}; // @[Cat.scala 29:58]
  assign _T_19 = $signed(_T_14) < 13'sh402; // @[fNFromRecFN.scala 50:39]
  assign _T_22 = 6'h1 - _T_14[5:0]; // @[fNFromRecFN.scala 51:39]
  assign _T_24 = _T_18[53:1] >> _T_22; // @[fNFromRecFN.scala 52:42]
  assign _T_28 = _T_14[10:0] - 11'h401; // @[fNFromRecFN.scala 57:45]
  assign _T_29 = _T_19 ? 11'h0 : _T_28; // @[fNFromRecFN.scala 55:16]
  assign _T_30 = _T_9 | _T_12; // @[fNFromRecFN.scala 59:44]
  assign _T_32 = _T_30 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  assign _T_33 = _T_29 | _T_32; // @[fNFromRecFN.scala 59:15]
  assign _T_35 = _T_12 ? 52'h0 : _T_18[51:0]; // @[fNFromRecFN.scala 63:20]
  assign _T_36 = _T_19 ? _T_24[51:0] : _T_35; // @[fNFromRecFN.scala 61:16]
  assign _T_38 = {in_in1[64],_T_33,_T_36}; // @[Cat.scala 29:58]
  assign _T_43 = {in_in1[31],in_in1[52],in_in1[30:0]}; // @[Cat.scala 29:58]
  assign _T_46 = _T_43[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_48 = _T_43[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign _T_51 = _T_48 & _T_43[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign _T_54 = _T_48 & ~_T_43[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign _T_56 = {1'b0,$signed(_T_43[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign _T_60 = {1'h0,~_T_46,_T_43[22:0]}; // @[Cat.scala 29:58]
  assign _T_61 = $signed(_T_56) < 10'sh82; // @[fNFromRecFN.scala 50:39]
  assign _T_64 = 5'h1 - _T_56[4:0]; // @[fNFromRecFN.scala 51:39]
  assign _T_66 = _T_60[24:1] >> _T_64; // @[fNFromRecFN.scala 52:42]
  assign _T_70 = _T_56[7:0] - 8'h81; // @[fNFromRecFN.scala 57:45]
  assign _T_71 = _T_61 ? 8'h0 : _T_70; // @[fNFromRecFN.scala 55:16]
  assign _T_72 = _T_51 | _T_54; // @[fNFromRecFN.scala 59:44]
  assign _T_74 = _T_72 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_75 = _T_71 | _T_74; // @[fNFromRecFN.scala 59:15]
  assign _T_77 = _T_54 ? 23'h0 : _T_60[22:0]; // @[fNFromRecFN.scala 63:20]
  assign _T_78 = _T_61 ? _T_66[22:0] : _T_77; // @[fNFromRecFN.scala 61:16]
  assign _T_80 = {_T_43[32],_T_75,_T_78}; // @[Cat.scala 29:58]
  assign _T_83 = &in_in1[63:61]; // @[FPU.scala 203:56]
  assign _T_85 = _T_83 ? _T_80 : _T_38[31:0]; // @[FPU.scala 394:44]
  assign store = {_T_38[63:32],_T_85}; // @[Cat.scala 29:58]
  assign _T_87 = {store[31:0],store[31:0]}; // @[Cat.scala 29:58]
  assign _T_247 = RecFNToIN_io_intExceptionFlags[2] | RecFNToIN_1_io_intExceptionFlags[1]; // @[FPU.scala 462:54]
  assign _T_239 = in_in1[64] & ~_T_83; // @[FPU.scala 460:59]
  assign _T_240 = RecFNToIN_io_signedOut == _T_239; // @[FPU.scala 461:46]
  assign _T_243 = _T_239 ? 31'h0 : 31'h7fffffff; // @[Bitwise.scala 72:12]
  assign _T_249 = {RecFNToIN_io_out[63:32],_T_240,_T_243}; // @[Cat.scala 29:58]
  assign _GEN_24 = _T_247 ? _T_249 : RecFNToIN_io_out; // @[FPU.scala 463:26]
  assign _GEN_25 = in_typ[1] ? RecFNToIN_io_out : _GEN_24; // @[FPU.scala 454:30]
  assign _T_217 = {dcmp_io_lt,dcmp_io_eq}; // @[Cat.scala 29:58]
  assign _GEN_33 = {{1'd0}, _T_217}; // @[FPU.scala 438:22]
  assign _T_218 = ~in_rm & _GEN_33; // @[FPU.scala 438:22]
  assign _T_219 = |_T_218; // @[FPU.scala 438:53]
  assign _T_221 = {store[63:32], 32'h0}; // @[FPU.scala 438:77]
  assign _GEN_34 = {{63'd0}, _T_219}; // @[FPU.scala 438:57]
  assign _T_222 = _GEN_34 | _T_221; // @[FPU.scala 438:57]
  assign _GEN_28 = in_ren2 ? _T_222 : _GEN_25; // @[FPU.scala 442:21]
  assign _T_189 = _T_83 & in_in1[51]; // @[FPU.scala 219:24]
  assign _T_187 = _T_83 & ~in_in1[51]; // @[FPU.scala 218:24]
  assign _T_168 = in_in1[63:62] == 2'h3; // @[FPU.scala 210:28]
  assign _T_183 = _T_168 & ~in_in1[61]; // @[FPU.scala 216:27]
  assign _T_191 = _T_183 & ~in_in1[64]; // @[FPU.scala 221:31]
  assign _T_175 = in_in1[63:62] == 2'h1; // @[FPU.scala 214:27]
  assign _T_170 = in_in1[61:52] < 10'h2; // @[FPU.scala 212:55]
  assign _T_177 = _T_175 & ~_T_170; // @[FPU.scala 214:39]
  assign _T_178 = in_in1[63:62] == 2'h2; // @[FPU.scala 214:71]
  assign _T_179 = _T_177 | _T_178; // @[FPU.scala 214:61]
  assign _T_193 = _T_179 & ~in_in1[64]; // @[FPU.scala 221:50]
  assign _T_171 = in_in1[63:61] == 3'h1; // @[FPU.scala 213:28]
  assign _T_173 = _T_175 & _T_170; // @[FPU.scala 213:62]
  assign _T_174 = _T_171 | _T_173; // @[FPU.scala 213:40]
  assign _T_195 = _T_174 & ~in_in1[64]; // @[FPU.scala 222:21]
  assign _T_180 = in_in1[63:61] == 3'h0; // @[FPU.scala 215:23]
  assign _T_197 = _T_180 & ~in_in1[64]; // @[FPU.scala 222:38]
  assign _T_198 = _T_180 & in_in1[64]; // @[FPU.scala 222:55]
  assign _T_199 = _T_174 & in_in1[64]; // @[FPU.scala 223:21]
  assign _T_200 = _T_179 & in_in1[64]; // @[FPU.scala 223:39]
  assign _T_201 = _T_183 & in_in1[64]; // @[FPU.scala 223:54]
  assign _T_210 = {_T_189,_T_187,_T_191,_T_193,_T_195,_T_197,_T_198,_T_199,_T_200,_T_201}; // @[Cat.scala 29:58]
  assign _T_111 = in_in1[63:61] >= 3'h6; // @[FPU.scala 235:36]
  assign _T_112 = _T_4 | _T_111; // @[FPU.scala 235:25]
  assign _T_107 = in_in1[63:52] + 12'h100; // @[FPU.scala 234:31]
  assign _T_109 = _T_107 - 12'h800; // @[FPU.scala 234:48]
  assign _T_114 = {in_in1[63:61],_T_109[5:0]}; // @[Cat.scala 29:58]
  assign _T_116 = _T_112 ? _T_114 : _T_109[8:0]; // @[FPU.scala 235:10]
  assign _T_103 = {in_in1[51:0], 24'h0}; // @[FPU.scala 231:28]
  assign _T_118 = {in_in1[64],_T_116,_T_103[75:53]}; // @[Cat.scala 29:58]
  assign _T_138 = &_T_118[31:29]; // @[FPU.scala 217:22]
  assign _T_143 = _T_138 & _T_118[22]; // @[FPU.scala 219:24]
  assign _T_141 = _T_138 & ~_T_118[22]; // @[FPU.scala 218:24]
  assign _T_122 = _T_118[31:30] == 2'h3; // @[FPU.scala 210:28]
  assign _T_137 = _T_122 & ~_T_118[29]; // @[FPU.scala 216:27]
  assign _T_145 = _T_137 & ~_T_118[32]; // @[FPU.scala 221:31]
  assign _T_129 = _T_118[31:30] == 2'h1; // @[FPU.scala 214:27]
  assign _T_124 = _T_118[29:23] < 7'h2; // @[FPU.scala 212:55]
  assign _T_131 = _T_129 & ~_T_124; // @[FPU.scala 214:39]
  assign _T_132 = _T_118[31:30] == 2'h2; // @[FPU.scala 214:71]
  assign _T_133 = _T_131 | _T_132; // @[FPU.scala 214:61]
  assign _T_147 = _T_133 & ~_T_118[32]; // @[FPU.scala 221:50]
  assign _T_125 = _T_118[31:29] == 3'h1; // @[FPU.scala 213:28]
  assign _T_127 = _T_129 & _T_124; // @[FPU.scala 213:62]
  assign _T_128 = _T_125 | _T_127; // @[FPU.scala 213:40]
  assign _T_149 = _T_128 & ~_T_118[32]; // @[FPU.scala 222:21]
  assign _T_134 = _T_118[31:29] == 3'h0; // @[FPU.scala 215:23]
  assign _T_151 = _T_134 & ~_T_118[32]; // @[FPU.scala 222:38]
  assign _T_152 = _T_134 & _T_118[32]; // @[FPU.scala 222:55]
  assign _T_153 = _T_128 & _T_118[32]; // @[FPU.scala 223:21]
  assign _T_154 = _T_133 & _T_118[32]; // @[FPU.scala 223:39]
  assign _T_155 = _T_137 & _T_118[32]; // @[FPU.scala 223:54]
  assign _T_164 = {_T_143,_T_141,_T_145,_T_147,_T_149,_T_151,_T_152,_T_153,_T_154,_T_155}; // @[Cat.scala 29:58]
  assign _T_212 = tag ? _T_210 : _T_164; // @[package.scala 32:76]
  assign _GEN_35 = {{54'd0}, _T_212}; // @[FPU.scala 433:27]
  assign _T_215 = _GEN_35 | _T_221; // @[FPU.scala 433:27]
  assign _GEN_22 = in_rm[0] ? _T_215 : store; // @[FPU.scala 431:19]
  assign toint = in_wflags ? _GEN_28 : _GEN_22; // @[FPU.scala 437:20]
  assign _T_94 = toint[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _T_95 = {_T_94,toint[31:0]}; // @[Cat.scala 29:58]
  assign _GEN_27 = ~in_ren2 & in_typ[1]; // @[FPU.scala 442:21]
  assign _GEN_23 = in_rm[0] ? 1'h0 : tag; // @[FPU.scala 431:19]
  assign intType = in_wflags ? _GEN_27 : _GEN_23; // @[FPU.scala 437:20]
  assign _T_228 = |RecFNToIN_io_intExceptionFlags[2:1]; // @[FPU.scala 450:62]
  assign _T_231 = {_T_228,3'h0,RecFNToIN_io_intExceptionFlags[0]}; // @[Cat.scala 29:58]
  assign _T_252 = ~_T_247 & RecFNToIN_io_intExceptionFlags[0]; // @[FPU.scala 464:64]
  assign _T_254 = {_T_247,3'h0,_T_252}; // @[Cat.scala 29:58]
  assign _GEN_26 = in_typ[1] ? _T_231 : _T_254; // @[FPU.scala 454:30]
  assign _GEN_29 = in_ren2 ? dcmp_io_exceptionFlags : _GEN_26; // @[FPU.scala 442:21]
  assign _T_256 = $signed(dcmp_io_a) < 65'sh0; // @[FPU.scala 471:53]
  assign _T_258 = $signed(dcmp_io_b) >= 65'sh0; // @[FPU.scala 471:79]
  assign _T_259 = _T_256 & _T_258; // @[FPU.scala 471:59]
  assign io_out_bits_in_rm = in_rm; // @[FPU.scala 472:18]
  assign io_out_bits_in_in1 = in_in1; // @[FPU.scala 472:18]
  assign io_out_bits_in_in2 = in_in2; // @[FPU.scala 472:18]
  assign io_out_bits_lt = dcmp_io_lt | _T_259; // @[FPU.scala 471:18]
  assign io_out_bits_store = tag ? store : _T_87; // @[FPU.scala 427:21]
  assign io_out_bits_toint = intType ? toint : _T_95; // @[FPU.scala 428:21]
  assign io_out_bits_exc = in_wflags ? _GEN_29 : 5'h0; // @[FPU.scala 429:19 FPU.scala 439:21 FPU.scala 450:23 FPU.scala 464:27]
  assign dcmp_io_a = in_in1; // @[FPU.scala 419:13]
  assign dcmp_io_b = in_in2; // @[FPU.scala 420:13]
  assign dcmp_io_signaling = ~in_rm[1]; // @[FPU.scala 421:21]
  assign RecFNToIN_io_in = in_in1; // @[FPU.scala 446:18]
  assign RecFNToIN_io_roundingMode = in_rm; // @[FPU.scala 447:28]
  assign RecFNToIN_io_signedOut = ~in_typ[0]; // @[FPU.scala 448:25]
  assign RecFNToIN_1_io_in = in_in1; // @[FPU.scala 456:24]
  assign RecFNToIN_1_io_roundingMode = in_rm; // @[FPU.scala 457:34]
  assign RecFNToIN_1_io_signedOut = ~in_typ[0]; // @[FPU.scala 458:31]
  assign FPToInt_cov_read_addr = FPToInt_state;
  assign FPToInt_cov_read_data = FPToInt_cov[FPToInt_cov_read_addr]; // @[Coverage map for FPToInt]
  assign FPToInt_cov_write_data = 1'h1;
  assign FPToInt_cov_write_addr = FPToInt_state;
  assign FPToInt_cov_write_mask = 1'h1;
  assign FPToInt_cov_write_en = 1'h1;
  assign in_wflags_shl = in_wflags;
  assign in_wflags_pad = {4'h0,in_wflags_shl};
  assign in_singleOut_shl = {in_singleOut, 1'h0};
  assign in_singleOut_pad = {3'h0,in_singleOut_shl};
  assign in_typ_shl = {in_typ, 2'h0};
  assign in_typ_pad = {1'h0,in_typ_shl};
  assign in_ren2_shl = {in_ren2, 4'h0};
  assign in_ren2_pad = in_ren2_shl;
  assign FPToInt_xor1 = in_wflags_pad ^ in_singleOut_pad;
  assign FPToInt_xor2 = in_typ_pad ^ in_ren2_pad;
  assign FPToInt_xor0 = FPToInt_xor1 ^ FPToInt_xor2;
  assign dcmp_sum = FPToInt_covSum + dcmp_io_covSum;
  assign RecFNToIN_sum = dcmp_sum + RecFNToIN_io_covSum;
  assign RecFNToIN_1_sum = RecFNToIN_sum + RecFNToIN_1_io_covSum;
  assign io_covSum = RecFNToIN_1_sum;
  assign dcmp_metaAssert_wire = dcmp_metaAssert;
  assign RecFNToIN_metaAssert_wire = RecFNToIN_metaAssert;
  assign RecFNToIN_1_metaAssert_wire = RecFNToIN_1_metaAssert;
  assign FPToInt_or2 = RecFNToIN_metaAssert_wire | RecFNToIN_1_metaAssert_wire;
  assign FPToInt_or0 = dcmp_metaAssert_wire | FPToInt_or2;
  assign metaAssert = FPToInt_or0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_ren2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_singleOut = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_wflags = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_rm = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_typ = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  in_in1 = _RAND_5[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  in_in2 = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  FPToInt_state = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    FPToInt_cov[initvar] = _RAND_8[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  FPToInt_covSum = _RAND_9[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      in_ren2 <= 1'h0;
    end else if (io_in_valid) begin
      in_ren2 <= io_in_bits_ren2;
    end
    if (metaReset) begin
      in_singleOut <= 1'h0;
    end else if (io_in_valid) begin
      in_singleOut <= io_in_bits_singleOut;
    end
    if (metaReset) begin
      in_wflags <= 1'h0;
    end else if (io_in_valid) begin
      in_wflags <= io_in_bits_wflags;
    end
    if (metaReset) begin
      in_rm <= 3'h0;
    end else if (io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      in_typ <= 2'h0;
    end else if (io_in_valid) begin
      in_typ <= io_in_bits_typ;
    end
    if (metaReset) begin
      in_in1 <= 65'h0;
    end else if (io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      in_in2 <= 65'h0;
    end else if (io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    FPToInt_state <= FPToInt_xor0;
    if (!(FPToInt_cov_read_data)) begin
      FPToInt_covSum <= FPToInt_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(FPToInt_cov_write_en & FPToInt_cov_write_mask) begin
      FPToInt_cov[FPToInt_cov_write_addr] <= FPToInt_cov_write_data; // @[Coverage map for FPToInt]
    end
  end
endmodule
module IntToFP(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_singleIn,
  input         io_in_bits_wflags,
  input  [2:0]  io_in_bits_rm,
  input  [1:0]  io_in_bits_typ,
  input  [63:0] io_in_bits_in1,
  output [64:0] io_out_bits_data,
  output [4:0]  io_out_bits_exc,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire  INToRecFN_io_signedIn; // @[FPU.scala 503:23]
  wire [63:0] INToRecFN_io_in; // @[FPU.scala 503:23]
  wire [2:0] INToRecFN_io_roundingMode; // @[FPU.scala 503:23]
  wire [32:0] INToRecFN_io_out; // @[FPU.scala 503:23]
  wire [4:0] INToRecFN_io_exceptionFlags; // @[FPU.scala 503:23]
  wire [29:0] INToRecFN_io_covSum; // @[FPU.scala 503:23]
  wire  INToRecFN_metaAssert; // @[FPU.scala 503:23]
  wire  INToRecFN_1_io_signedIn; // @[FPU.scala 503:23]
  wire [63:0] INToRecFN_1_io_in; // @[FPU.scala 503:23]
  wire [2:0] INToRecFN_1_io_roundingMode; // @[FPU.scala 503:23]
  wire [64:0] INToRecFN_1_io_out; // @[FPU.scala 503:23]
  wire [4:0] INToRecFN_1_io_exceptionFlags; // @[FPU.scala 503:23]
  wire [29:0] INToRecFN_1_io_covSum; // @[FPU.scala 503:23]
  wire  INToRecFN_1_metaAssert; // @[FPU.scala 503:23]
  reg  inPipe_valid; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg  inPipe_bits_singleIn; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  inPipe_bits_wflags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [2:0] inPipe_bits_rm; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [1:0] inPipe_bits_typ; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [63:0] inPipe_bits_in1; // @[Reg.scala 15:16]
  reg [63:0] _RAND_5;
  wire  tag; // @[FPU.scala 482:13]
  wire [63:0] _T_2; // @[package.scala 32:76]
  wire [63:0] _T_3; // @[FPU.scala 379:23]
  wire  _T_7; // @[rawFloatFromFN.scala 50:34]
  wire  _T_8; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_61; // @[Mux.scala 47:69]
  wire [5:0] _T_62; // @[Mux.scala 47:69]
  wire [5:0] _T_63; // @[Mux.scala 47:69]
  wire [5:0] _T_64; // @[Mux.scala 47:69]
  wire [5:0] _T_65; // @[Mux.scala 47:69]
  wire [5:0] _T_66; // @[Mux.scala 47:69]
  wire [5:0] _T_67; // @[Mux.scala 47:69]
  wire [5:0] _T_68; // @[Mux.scala 47:69]
  wire [5:0] _T_69; // @[Mux.scala 47:69]
  wire [5:0] _T_70; // @[Mux.scala 47:69]
  wire [5:0] _T_71; // @[Mux.scala 47:69]
  wire [5:0] _T_72; // @[Mux.scala 47:69]
  wire [5:0] _T_73; // @[Mux.scala 47:69]
  wire [5:0] _T_74; // @[Mux.scala 47:69]
  wire [5:0] _T_75; // @[Mux.scala 47:69]
  wire [5:0] _T_76; // @[Mux.scala 47:69]
  wire [5:0] _T_77; // @[Mux.scala 47:69]
  wire [5:0] _T_78; // @[Mux.scala 47:69]
  wire [5:0] _T_79; // @[Mux.scala 47:69]
  wire [5:0] _T_80; // @[Mux.scala 47:69]
  wire [5:0] _T_81; // @[Mux.scala 47:69]
  wire [5:0] _T_82; // @[Mux.scala 47:69]
  wire [5:0] _T_83; // @[Mux.scala 47:69]
  wire [5:0] _T_84; // @[Mux.scala 47:69]
  wire [5:0] _T_85; // @[Mux.scala 47:69]
  wire [5:0] _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_106; // @[Mux.scala 47:69]
  wire [5:0] _T_107; // @[Mux.scala 47:69]
  wire [5:0] _T_108; // @[Mux.scala 47:69]
  wire [5:0] _T_109; // @[Mux.scala 47:69]
  wire [5:0] _T_110; // @[Mux.scala 47:69]
  wire [5:0] _T_111; // @[Mux.scala 47:69]
  wire [114:0] _GEN_24; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_112; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_114; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_25; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_115; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_116; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_117; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_26; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_118; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_27; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_120; // @[rawFloatFromFN.scala 59:15]
  wire  _T_121; // @[rawFloatFromFN.scala 62:34]
  wire  _T_123; // @[rawFloatFromFN.scala 63:62]
  wire  _T_126; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_129; // @[rawFloatFromFN.scala 70:48]
  wire [51:0] _T_131; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_133; // @[Cat.scala 29:58]
  wire [2:0] _T_135; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_28; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_137; // @[recFNFromFN.scala 48:79]
  wire [64:0] _T_142; // @[Cat.scala 29:58]
  wire  _T_146; // @[rawFloatFromFN.scala 50:34]
  wire  _T_147; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_171; // @[Mux.scala 47:69]
  wire [4:0] _T_172; // @[Mux.scala 47:69]
  wire [4:0] _T_173; // @[Mux.scala 47:69]
  wire [4:0] _T_174; // @[Mux.scala 47:69]
  wire [4:0] _T_175; // @[Mux.scala 47:69]
  wire [4:0] _T_176; // @[Mux.scala 47:69]
  wire [4:0] _T_177; // @[Mux.scala 47:69]
  wire [4:0] _T_178; // @[Mux.scala 47:69]
  wire [4:0] _T_179; // @[Mux.scala 47:69]
  wire [4:0] _T_180; // @[Mux.scala 47:69]
  wire [4:0] _T_181; // @[Mux.scala 47:69]
  wire [4:0] _T_182; // @[Mux.scala 47:69]
  wire [4:0] _T_183; // @[Mux.scala 47:69]
  wire [4:0] _T_184; // @[Mux.scala 47:69]
  wire [4:0] _T_185; // @[Mux.scala 47:69]
  wire [4:0] _T_186; // @[Mux.scala 47:69]
  wire [4:0] _T_187; // @[Mux.scala 47:69]
  wire [4:0] _T_188; // @[Mux.scala 47:69]
  wire [4:0] _T_189; // @[Mux.scala 47:69]
  wire [4:0] _T_190; // @[Mux.scala 47:69]
  wire [4:0] _T_191; // @[Mux.scala 47:69]
  wire [4:0] _T_192; // @[Mux.scala 47:69]
  wire [53:0] _GEN_29; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_193; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_195; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_30; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_196; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_197; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_198; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_31; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_199; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_32; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_201; // @[rawFloatFromFN.scala 59:15]
  wire  _T_202; // @[rawFloatFromFN.scala 62:34]
  wire  _T_204; // @[rawFloatFromFN.scala 63:62]
  wire  _T_207; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_210; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_212; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_214; // @[Cat.scala 29:58]
  wire [2:0] _T_216; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_33; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_218; // @[recFNFromFN.scala 48:79]
  wire [32:0] _T_223; // @[Cat.scala 29:58]
  wire  _T_226; // @[FPU.scala 286:42]
  wire [64:0] _T_237; // @[Cat.scala 29:58]
  wire  _T_239; // @[FPU.scala 203:56]
  wire [32:0] _T_247; // @[FPU.scala 493:45]
  wire [31:0] _T_248; // @[FPU.scala 493:60]
  wire [32:0] _T_249; // @[FPU.scala 493:19]
  wire [64:0] _T_255; // @[FPU.scala 361:25]
  wire  _T_257; // @[FPU.scala 203:56]
  wire [64:0] _T_258; // @[FPU.scala 362:10]
  wire [64:0] _T_260; // @[Cat.scala 29:58]
  reg [64:0] _T_266_data; // @[Reg.scala 15:16]
  reg [95:0] _RAND_6;
  reg [4:0] _T_266_exc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [4:0] IntToFP_state; // @[Register tracking IntToFP state]
  reg [31:0] _RAND_8;
  reg  IntToFP_cov [0:31]; // @[Coverage map for IntToFP]
  reg [31:0] _RAND_9;
  wire  IntToFP_cov_read_data; // @[Coverage map for IntToFP]
  wire [4:0] IntToFP_cov_read_addr; // @[Coverage map for IntToFP]
  wire  IntToFP_cov_write_data; // @[Coverage map for IntToFP]
  wire [4:0] IntToFP_cov_write_addr; // @[Coverage map for IntToFP]
  wire  IntToFP_cov_write_mask; // @[Coverage map for IntToFP]
  wire  IntToFP_cov_write_en; // @[Coverage map for IntToFP]
  reg [29:0] IntToFP_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_10;
  wire  inPipe_bits_singleIn_shl;
  wire [4:0] inPipe_bits_singleIn_pad;
  wire [1:0] inPipe_valid_shl;
  wire [4:0] inPipe_valid_pad;
  wire [2:0] inPipe_bits_wflags_shl;
  wire [4:0] inPipe_bits_wflags_pad;
  wire [4:0] inPipe_bits_typ_shl;
  wire [4:0] inPipe_bits_typ_pad;
  wire [4:0] IntToFP_xor1;
  wire [4:0] IntToFP_xor2;
  wire [4:0] IntToFP_xor0;
  wire [29:0] INToRecFN_sum;
  wire [29:0] INToRecFN_1_sum;
  wire  INToRecFN_metaAssert_wire;
  wire  INToRecFN_1_metaAssert_wire;
  wire  IntToFP_or0;
  reg  IntToFP_metaAssert;
  reg [31:0] _RAND_11;
  INToRecFN INToRecFN ( // @[FPU.scala 503:23]
    .io_signedIn(INToRecFN_io_signedIn),
    .io_in(INToRecFN_io_in),
    .io_roundingMode(INToRecFN_io_roundingMode),
    .io_out(INToRecFN_io_out),
    .io_exceptionFlags(INToRecFN_io_exceptionFlags),
    .io_covSum(INToRecFN_io_covSum),
    .metaAssert(INToRecFN_metaAssert)
  );
  INToRecFN_1 INToRecFN_1 ( // @[FPU.scala 503:23]
    .io_signedIn(INToRecFN_1_io_signedIn),
    .io_in(INToRecFN_1_io_in),
    .io_roundingMode(INToRecFN_1_io_roundingMode),
    .io_out(INToRecFN_1_io_out),
    .io_exceptionFlags(INToRecFN_1_io_exceptionFlags),
    .io_covSum(INToRecFN_1_io_covSum),
    .metaAssert(INToRecFN_1_metaAssert)
  );
  assign tag = ~inPipe_bits_singleIn; // @[FPU.scala 482:13]
  assign _T_2 = tag ? 64'h0 : 64'hffffffff00000000; // @[package.scala 32:76]
  assign _T_3 = _T_2 | inPipe_bits_in1; // @[FPU.scala 379:23]
  assign _T_7 = _T_3[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_8 = _T_3[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_61 = _T_3[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  assign _T_62 = _T_3[2] ? 6'h31 : _T_61; // @[Mux.scala 47:69]
  assign _T_63 = _T_3[3] ? 6'h30 : _T_62; // @[Mux.scala 47:69]
  assign _T_64 = _T_3[4] ? 6'h2f : _T_63; // @[Mux.scala 47:69]
  assign _T_65 = _T_3[5] ? 6'h2e : _T_64; // @[Mux.scala 47:69]
  assign _T_66 = _T_3[6] ? 6'h2d : _T_65; // @[Mux.scala 47:69]
  assign _T_67 = _T_3[7] ? 6'h2c : _T_66; // @[Mux.scala 47:69]
  assign _T_68 = _T_3[8] ? 6'h2b : _T_67; // @[Mux.scala 47:69]
  assign _T_69 = _T_3[9] ? 6'h2a : _T_68; // @[Mux.scala 47:69]
  assign _T_70 = _T_3[10] ? 6'h29 : _T_69; // @[Mux.scala 47:69]
  assign _T_71 = _T_3[11] ? 6'h28 : _T_70; // @[Mux.scala 47:69]
  assign _T_72 = _T_3[12] ? 6'h27 : _T_71; // @[Mux.scala 47:69]
  assign _T_73 = _T_3[13] ? 6'h26 : _T_72; // @[Mux.scala 47:69]
  assign _T_74 = _T_3[14] ? 6'h25 : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = _T_3[15] ? 6'h24 : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = _T_3[16] ? 6'h23 : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = _T_3[17] ? 6'h22 : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = _T_3[18] ? 6'h21 : _T_77; // @[Mux.scala 47:69]
  assign _T_79 = _T_3[19] ? 6'h20 : _T_78; // @[Mux.scala 47:69]
  assign _T_80 = _T_3[20] ? 6'h1f : _T_79; // @[Mux.scala 47:69]
  assign _T_81 = _T_3[21] ? 6'h1e : _T_80; // @[Mux.scala 47:69]
  assign _T_82 = _T_3[22] ? 6'h1d : _T_81; // @[Mux.scala 47:69]
  assign _T_83 = _T_3[23] ? 6'h1c : _T_82; // @[Mux.scala 47:69]
  assign _T_84 = _T_3[24] ? 6'h1b : _T_83; // @[Mux.scala 47:69]
  assign _T_85 = _T_3[25] ? 6'h1a : _T_84; // @[Mux.scala 47:69]
  assign _T_86 = _T_3[26] ? 6'h19 : _T_85; // @[Mux.scala 47:69]
  assign _T_87 = _T_3[27] ? 6'h18 : _T_86; // @[Mux.scala 47:69]
  assign _T_88 = _T_3[28] ? 6'h17 : _T_87; // @[Mux.scala 47:69]
  assign _T_89 = _T_3[29] ? 6'h16 : _T_88; // @[Mux.scala 47:69]
  assign _T_90 = _T_3[30] ? 6'h15 : _T_89; // @[Mux.scala 47:69]
  assign _T_91 = _T_3[31] ? 6'h14 : _T_90; // @[Mux.scala 47:69]
  assign _T_92 = _T_3[32] ? 6'h13 : _T_91; // @[Mux.scala 47:69]
  assign _T_93 = _T_3[33] ? 6'h12 : _T_92; // @[Mux.scala 47:69]
  assign _T_94 = _T_3[34] ? 6'h11 : _T_93; // @[Mux.scala 47:69]
  assign _T_95 = _T_3[35] ? 6'h10 : _T_94; // @[Mux.scala 47:69]
  assign _T_96 = _T_3[36] ? 6'hf : _T_95; // @[Mux.scala 47:69]
  assign _T_97 = _T_3[37] ? 6'he : _T_96; // @[Mux.scala 47:69]
  assign _T_98 = _T_3[38] ? 6'hd : _T_97; // @[Mux.scala 47:69]
  assign _T_99 = _T_3[39] ? 6'hc : _T_98; // @[Mux.scala 47:69]
  assign _T_100 = _T_3[40] ? 6'hb : _T_99; // @[Mux.scala 47:69]
  assign _T_101 = _T_3[41] ? 6'ha : _T_100; // @[Mux.scala 47:69]
  assign _T_102 = _T_3[42] ? 6'h9 : _T_101; // @[Mux.scala 47:69]
  assign _T_103 = _T_3[43] ? 6'h8 : _T_102; // @[Mux.scala 47:69]
  assign _T_104 = _T_3[44] ? 6'h7 : _T_103; // @[Mux.scala 47:69]
  assign _T_105 = _T_3[45] ? 6'h6 : _T_104; // @[Mux.scala 47:69]
  assign _T_106 = _T_3[46] ? 6'h5 : _T_105; // @[Mux.scala 47:69]
  assign _T_107 = _T_3[47] ? 6'h4 : _T_106; // @[Mux.scala 47:69]
  assign _T_108 = _T_3[48] ? 6'h3 : _T_107; // @[Mux.scala 47:69]
  assign _T_109 = _T_3[49] ? 6'h2 : _T_108; // @[Mux.scala 47:69]
  assign _T_110 = _T_3[50] ? 6'h1 : _T_109; // @[Mux.scala 47:69]
  assign _T_111 = _T_3[51] ? 6'h0 : _T_110; // @[Mux.scala 47:69]
  assign _GEN_24 = {{63'd0}, _T_3[51:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_112 = _GEN_24 << _T_111; // @[rawFloatFromFN.scala 54:36]
  assign _T_114 = {_T_112[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_25 = {{6'd0}, _T_111}; // @[rawFloatFromFN.scala 57:26]
  assign _T_115 = _GEN_25 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _T_116 = _T_7 ? _T_115 : {{1'd0}, _T_3[62:52]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_117 = _T_7 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_26 = {{9'd0}, _T_117}; // @[rawFloatFromFN.scala 60:22]
  assign _T_118 = 11'h400 | _GEN_26; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_27 = {{1'd0}, _T_118}; // @[rawFloatFromFN.scala 59:15]
  assign _T_120 = _T_116 + _GEN_27; // @[rawFloatFromFN.scala 59:15]
  assign _T_121 = _T_7 & _T_8; // @[rawFloatFromFN.scala 62:34]
  assign _T_123 = _T_120[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_126 = _T_123 & ~_T_8; // @[rawFloatFromFN.scala 66:33]
  assign _T_129 = {1'b0,$signed(_T_120)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_131 = _T_7 ? _T_114 : _T_3[51:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_133 = {1'h0,~_T_121,_T_131}; // @[Cat.scala 29:58]
  assign _T_135 = _T_121 ? 3'h0 : _T_129[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_28 = {{2'd0}, _T_126}; // @[recFNFromFN.scala 48:79]
  assign _T_137 = _T_135 | _GEN_28; // @[recFNFromFN.scala 48:79]
  assign _T_142 = {_T_3[63],_T_137,_T_129[8:0],_T_133[51:0]}; // @[Cat.scala 29:58]
  assign _T_146 = _T_3[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_147 = _T_3[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_171 = _T_3[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _T_172 = _T_3[2] ? 5'h14 : _T_171; // @[Mux.scala 47:69]
  assign _T_173 = _T_3[3] ? 5'h13 : _T_172; // @[Mux.scala 47:69]
  assign _T_174 = _T_3[4] ? 5'h12 : _T_173; // @[Mux.scala 47:69]
  assign _T_175 = _T_3[5] ? 5'h11 : _T_174; // @[Mux.scala 47:69]
  assign _T_176 = _T_3[6] ? 5'h10 : _T_175; // @[Mux.scala 47:69]
  assign _T_177 = _T_3[7] ? 5'hf : _T_176; // @[Mux.scala 47:69]
  assign _T_178 = _T_3[8] ? 5'he : _T_177; // @[Mux.scala 47:69]
  assign _T_179 = _T_3[9] ? 5'hd : _T_178; // @[Mux.scala 47:69]
  assign _T_180 = _T_3[10] ? 5'hc : _T_179; // @[Mux.scala 47:69]
  assign _T_181 = _T_3[11] ? 5'hb : _T_180; // @[Mux.scala 47:69]
  assign _T_182 = _T_3[12] ? 5'ha : _T_181; // @[Mux.scala 47:69]
  assign _T_183 = _T_3[13] ? 5'h9 : _T_182; // @[Mux.scala 47:69]
  assign _T_184 = _T_3[14] ? 5'h8 : _T_183; // @[Mux.scala 47:69]
  assign _T_185 = _T_3[15] ? 5'h7 : _T_184; // @[Mux.scala 47:69]
  assign _T_186 = _T_3[16] ? 5'h6 : _T_185; // @[Mux.scala 47:69]
  assign _T_187 = _T_3[17] ? 5'h5 : _T_186; // @[Mux.scala 47:69]
  assign _T_188 = _T_3[18] ? 5'h4 : _T_187; // @[Mux.scala 47:69]
  assign _T_189 = _T_3[19] ? 5'h3 : _T_188; // @[Mux.scala 47:69]
  assign _T_190 = _T_3[20] ? 5'h2 : _T_189; // @[Mux.scala 47:69]
  assign _T_191 = _T_3[21] ? 5'h1 : _T_190; // @[Mux.scala 47:69]
  assign _T_192 = _T_3[22] ? 5'h0 : _T_191; // @[Mux.scala 47:69]
  assign _GEN_29 = {{31'd0}, _T_3[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_193 = _GEN_29 << _T_192; // @[rawFloatFromFN.scala 54:36]
  assign _T_195 = {_T_193[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_30 = {{4'd0}, _T_192}; // @[rawFloatFromFN.scala 57:26]
  assign _T_196 = _GEN_30 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_197 = _T_146 ? _T_196 : {{1'd0}, _T_3[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_198 = _T_146 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_31 = {{6'd0}, _T_198}; // @[rawFloatFromFN.scala 60:22]
  assign _T_199 = 8'h80 | _GEN_31; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_32 = {{1'd0}, _T_199}; // @[rawFloatFromFN.scala 59:15]
  assign _T_201 = _T_197 + _GEN_32; // @[rawFloatFromFN.scala 59:15]
  assign _T_202 = _T_146 & _T_147; // @[rawFloatFromFN.scala 62:34]
  assign _T_204 = _T_201[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_207 = _T_204 & ~_T_147; // @[rawFloatFromFN.scala 66:33]
  assign _T_210 = {1'b0,$signed(_T_201)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_212 = _T_146 ? _T_195 : _T_3[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_214 = {1'h0,~_T_202,_T_212}; // @[Cat.scala 29:58]
  assign _T_216 = _T_202 ? 3'h0 : _T_210[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_33 = {{2'd0}, _T_207}; // @[recFNFromFN.scala 48:79]
  assign _T_218 = _T_216 | _GEN_33; // @[recFNFromFN.scala 48:79]
  assign _T_223 = {_T_3[31],_T_218,_T_210[5:0],_T_214[22:0]}; // @[Cat.scala 29:58]
  assign _T_226 = &_T_142[51:32]; // @[FPU.scala 286:42]
  assign _T_237 = {_T_142[64:61],_T_226,_T_142[59:53],_T_223[31],_T_142[51:32],_T_223[32],_T_223[30:0]}; // @[Cat.scala 29:58]
  assign _T_239 = &_T_142[63:61]; // @[FPU.scala 203:56]
  assign _T_247 = {1'b0,$signed(inPipe_bits_in1[31:0])}; // @[FPU.scala 493:45]
  assign _T_248 = inPipe_bits_in1[31:0]; // @[FPU.scala 493:60]
  assign _T_249 = inPipe_bits_typ[0] ? $signed(_T_247) : $signed({{1{_T_248[31]}},_T_248}); // @[FPU.scala 493:19]
  assign _T_255 = INToRecFN_1_io_out & 65'h1efefffffffffffff; // @[FPU.scala 361:25]
  assign _T_257 = &INToRecFN_1_io_out[63:61]; // @[FPU.scala 203:56]
  assign _T_258 = _T_257 ? _T_255 : INToRecFN_1_io_out; // @[FPU.scala 362:10]
  assign _T_260 = {_T_258[64:33],INToRecFN_io_out}; // @[Cat.scala 29:58]
  assign io_out_bits_data = _T_266_data; // @[FPU.scala 517:10]
  assign io_out_bits_exc = _T_266_exc; // @[FPU.scala 517:10]
  assign INToRecFN_io_signedIn = ~inPipe_bits_typ[0]; // @[FPU.scala 504:23]
  assign INToRecFN_io_in = inPipe_bits_typ[1] ? $signed(inPipe_bits_in1) : $signed({{31{_T_249[32]}},_T_249}); // @[FPU.scala 505:17]
  assign INToRecFN_io_roundingMode = inPipe_bits_rm; // @[FPU.scala 506:27]
  assign INToRecFN_1_io_signedIn = ~inPipe_bits_typ[0]; // @[FPU.scala 504:23]
  assign INToRecFN_1_io_in = inPipe_bits_typ[1] ? $signed(inPipe_bits_in1) : $signed({{31{_T_249[32]}},_T_249}); // @[FPU.scala 505:17]
  assign INToRecFN_1_io_roundingMode = inPipe_bits_rm; // @[FPU.scala 506:27]
  assign IntToFP_cov_read_addr = IntToFP_state;
  assign IntToFP_cov_read_data = IntToFP_cov[IntToFP_cov_read_addr]; // @[Coverage map for IntToFP]
  assign IntToFP_cov_write_data = 1'h1;
  assign IntToFP_cov_write_addr = IntToFP_state;
  assign IntToFP_cov_write_mask = 1'h1;
  assign IntToFP_cov_write_en = 1'h1;
  assign inPipe_bits_singleIn_shl = inPipe_bits_singleIn;
  assign inPipe_bits_singleIn_pad = {4'h0,inPipe_bits_singleIn_shl};
  assign inPipe_valid_shl = {inPipe_valid, 1'h0};
  assign inPipe_valid_pad = {3'h0,inPipe_valid_shl};
  assign inPipe_bits_wflags_shl = {inPipe_bits_wflags, 2'h0};
  assign inPipe_bits_wflags_pad = {2'h0,inPipe_bits_wflags_shl};
  assign inPipe_bits_typ_shl = {inPipe_bits_typ, 3'h0};
  assign inPipe_bits_typ_pad = inPipe_bits_typ_shl;
  assign IntToFP_xor1 = inPipe_bits_singleIn_pad ^ inPipe_valid_pad;
  assign IntToFP_xor2 = inPipe_bits_wflags_pad ^ inPipe_bits_typ_pad;
  assign IntToFP_xor0 = IntToFP_xor1 ^ IntToFP_xor2;
  assign INToRecFN_sum = IntToFP_covSum + INToRecFN_io_covSum;
  assign INToRecFN_1_sum = INToRecFN_sum + INToRecFN_1_io_covSum;
  assign io_covSum = INToRecFN_1_sum;
  assign INToRecFN_metaAssert_wire = INToRecFN_metaAssert;
  assign INToRecFN_1_metaAssert_wire = INToRecFN_1_metaAssert;
  assign IntToFP_or0 = INToRecFN_metaAssert_wire | INToRecFN_1_metaAssert_wire;
  assign metaAssert = IntToFP_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inPipe_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inPipe_bits_singleIn = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  inPipe_bits_wflags = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  inPipe_bits_rm = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  inPipe_bits_typ = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  inPipe_bits_in1 = _RAND_5[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  _T_266_data = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_266_exc = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  IntToFP_state = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    IntToFP_cov[initvar] = _RAND_9[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  IntToFP_covSum = _RAND_10[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  IntToFP_metaAssert = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      inPipe_valid <= 1'h0;
    end else if (reset) begin
      inPipe_valid <= 1'h0;
    end else begin
      inPipe_valid <= io_in_valid;
    end
    if (metaReset) begin
      inPipe_bits_singleIn <= 1'h0;
    end else if (io_in_valid) begin
      inPipe_bits_singleIn <= io_in_bits_singleIn;
    end
    if (metaReset) begin
      inPipe_bits_wflags <= 1'h0;
    end else if (io_in_valid) begin
      inPipe_bits_wflags <= io_in_bits_wflags;
    end
    if (metaReset) begin
      inPipe_bits_rm <= 3'h0;
    end else if (io_in_valid) begin
      inPipe_bits_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      inPipe_bits_typ <= 2'h0;
    end else if (io_in_valid) begin
      inPipe_bits_typ <= io_in_bits_typ;
    end
    if (metaReset) begin
      inPipe_bits_in1 <= 64'h0;
    end else if (io_in_valid) begin
      inPipe_bits_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      _T_266_data <= 65'h0;
    end else if (inPipe_valid) begin
      if (inPipe_bits_wflags) begin
        if (tag) begin
          if (_T_257) begin
            _T_266_data <= _T_255;
          end else begin
            _T_266_data <= INToRecFN_1_io_out;
          end
        end else begin
          _T_266_data <= _T_260;
        end
      end else if (_T_239) begin
        _T_266_data <= _T_237;
      end else begin
        _T_266_data <= _T_142;
      end
    end
    if (metaReset) begin
      _T_266_exc <= 5'h0;
    end else if (inPipe_valid) begin
      if (inPipe_bits_wflags) begin
        if (tag) begin
          _T_266_exc <= INToRecFN_1_io_exceptionFlags;
        end else begin
          _T_266_exc <= INToRecFN_io_exceptionFlags;
        end
      end else begin
        _T_266_exc <= 5'h0;
      end
    end
    IntToFP_state <= IntToFP_xor0;
    if (!(IntToFP_cov_read_data)) begin
      IntToFP_covSum <= IntToFP_covSum + 1'h1;
    end
    if (metaReset) begin
      IntToFP_metaAssert <= 1'h0;
    end else begin
      IntToFP_metaAssert <= IntToFP_metaAssert | IntToFP_or0;
    end
  end
  always @(posedge clock) begin
    if(IntToFP_cov_write_en & IntToFP_cov_write_mask) begin
      IntToFP_cov[IntToFP_cov_write_addr] <= IntToFP_cov_write_data; // @[Coverage map for IntToFP]
    end
  end
endmodule
module FPToFP(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_ren2,
  input         io_in_bits_singleOut,
  input         io_in_bits_wflags,
  input  [2:0]  io_in_bits_rm,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  output [64:0] io_out_bits_data,
  output [4:0]  io_out_bits_exc,
  input         io_lt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [64:0] RecFNToRecFN_io_in; // @[FPU.scala 566:30]
  wire [2:0] RecFNToRecFN_io_roundingMode; // @[FPU.scala 566:30]
  wire [32:0] RecFNToRecFN_io_out; // @[FPU.scala 566:30]
  wire [4:0] RecFNToRecFN_io_exceptionFlags; // @[FPU.scala 566:30]
  wire [29:0] RecFNToRecFN_io_covSum; // @[FPU.scala 566:30]
  wire  RecFNToRecFN_metaAssert; // @[FPU.scala 566:30]
  reg  inPipe_valid; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg  inPipe_bits_ren2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  inPipe_bits_singleOut; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg  inPipe_bits_wflags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [2:0] inPipe_bits_rm; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [64:0] inPipe_bits_in1; // @[Reg.scala 15:16]
  reg [95:0] _RAND_5;
  reg [64:0] inPipe_bits_in2; // @[Reg.scala 15:16]
  reg [95:0] _RAND_6;
  wire [64:0] _T_1; // @[FPU.scala 529:48]
  wire [64:0] _T_4; // @[FPU.scala 529:66]
  wire [64:0] signNum; // @[FPU.scala 529:20]
  wire [64:0] fsgnj; // @[Cat.scala 29:58]
  wire  _T_8; // @[FPU.scala 203:56]
  wire  _T_10; // @[FPU.scala 203:56]
  wire  _T_15; // @[FPU.scala 204:34]
  wire  _T_20; // @[FPU.scala 204:34]
  wire  _T_21; // @[FPU.scala 539:49]
  wire  _T_22; // @[FPU.scala 540:27]
  wire  _T_24; // @[FPU.scala 541:41]
  wire  _T_26; // @[FPU.scala 541:51]
  wire  _T_27; // @[FPU.scala 541:24]
  wire [4:0] _T_28; // @[FPU.scala 542:31]
  wire [64:0] _T_29; // @[FPU.scala 543:53]
  wire [64:0] _T_30; // @[FPU.scala 543:25]
  wire [64:0] _GEN_23; // @[FPU.scala 536:25]
  wire  outTag; // @[FPU.scala 547:16]
  wire  _T_54; // @[FPU.scala 555:24]
  wire [64:0] _T_57; // @[FPU.scala 558:24]
  wire [64:0] fsgnjMux_data; // @[FPU.scala 555:42]
  wire [75:0] _T_36; // @[FPU.scala 231:28]
  wire [11:0] _T_40; // @[FPU.scala 234:31]
  wire [11:0] _T_42; // @[FPU.scala 234:48]
  wire  _T_43; // @[FPU.scala 235:19]
  wire  _T_44; // @[FPU.scala 235:36]
  wire  _T_45; // @[FPU.scala 235:25]
  wire [8:0] _T_47; // @[Cat.scala 29:58]
  wire [8:0] _T_49; // @[FPU.scala 235:10]
  wire [64:0] _T_52; // @[Cat.scala 29:58]
  wire [4:0] _T_63; // @[FPU.scala 560:51]
  wire [64:0] _T_69; // @[Cat.scala 29:58]
  reg [64:0] _T_71_data; // @[Reg.scala 15:16]
  reg [95:0] _RAND_7;
  reg [4:0] _T_71_exc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [6:0] FPToFP_state; // @[Register tracking FPToFP state]
  reg [31:0] _RAND_9;
  reg  FPToFP_cov [0:127]; // @[Coverage map for FPToFP]
  reg [31:0] _RAND_10;
  wire  FPToFP_cov_read_data; // @[Coverage map for FPToFP]
  wire [6:0] FPToFP_cov_read_addr; // @[Coverage map for FPToFP]
  wire  FPToFP_cov_write_data; // @[Coverage map for FPToFP]
  wire [6:0] FPToFP_cov_write_addr; // @[Coverage map for FPToFP]
  wire  FPToFP_cov_write_mask; // @[Coverage map for FPToFP]
  wire  FPToFP_cov_write_en; // @[Coverage map for FPToFP]
  reg [29:0] FPToFP_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_11;
  wire  inPipe_valid_shl;
  wire [6:0] inPipe_valid_pad;
  wire [1:0] inPipe_bits_singleOut_shl;
  wire [6:0] inPipe_bits_singleOut_pad;
  wire [2:0] inPipe_bits_ren2_shl;
  wire [6:0] inPipe_bits_ren2_pad;
  wire [3:0] inPipe_bits_wflags_shl;
  wire [6:0] inPipe_bits_wflags_pad;
  wire [6:0] inPipe_bits_rm_shl;
  wire [6:0] inPipe_bits_rm_pad;
  wire [6:0] FPToFP_xor1;
  wire [6:0] FPToFP_xor6;
  wire [6:0] FPToFP_xor2;
  wire [6:0] FPToFP_xor0;
  wire [29:0] RecFNToRecFN_sum;
  wire  RecFNToRecFN_metaAssert_wire;
  reg  FPToFP_metaAssert;
  reg [31:0] _RAND_12;
  RecFNToRecFN RecFNToRecFN ( // @[FPU.scala 566:30]
    .io_in(RecFNToRecFN_io_in),
    .io_roundingMode(RecFNToRecFN_io_roundingMode),
    .io_out(RecFNToRecFN_io_out),
    .io_exceptionFlags(RecFNToRecFN_io_exceptionFlags),
    .io_covSum(RecFNToRecFN_io_covSum),
    .metaAssert(RecFNToRecFN_metaAssert)
  );
  assign _T_1 = inPipe_bits_in1 ^ inPipe_bits_in2; // @[FPU.scala 529:48]
  assign _T_4 = inPipe_bits_rm[0] ? ~inPipe_bits_in2 : inPipe_bits_in2; // @[FPU.scala 529:66]
  assign signNum = inPipe_bits_rm[1] ? _T_1 : _T_4; // @[FPU.scala 529:20]
  assign fsgnj = {signNum[64],inPipe_bits_in1[63:0]}; // @[Cat.scala 29:58]
  assign _T_8 = &inPipe_bits_in1[63:61]; // @[FPU.scala 203:56]
  assign _T_10 = &inPipe_bits_in2[63:61]; // @[FPU.scala 203:56]
  assign _T_15 = _T_8 & ~inPipe_bits_in1[51]; // @[FPU.scala 204:34]
  assign _T_20 = _T_10 & ~inPipe_bits_in2[51]; // @[FPU.scala 204:34]
  assign _T_21 = _T_15 | _T_20; // @[FPU.scala 539:49]
  assign _T_22 = _T_8 & _T_10; // @[FPU.scala 540:27]
  assign _T_24 = inPipe_bits_rm[0] != io_lt; // @[FPU.scala 541:41]
  assign _T_26 = _T_24 & ~_T_8; // @[FPU.scala 541:51]
  assign _T_27 = _T_10 | _T_26; // @[FPU.scala 541:24]
  assign _T_28 = {_T_21, 4'h0}; // @[FPU.scala 542:31]
  assign _T_29 = _T_27 ? inPipe_bits_in1 : inPipe_bits_in2; // @[FPU.scala 543:53]
  assign _T_30 = _T_22 ? 65'he008000000000000 : _T_29; // @[FPU.scala 543:25]
  assign _GEN_23 = inPipe_bits_wflags ? _T_30 : fsgnj; // @[FPU.scala 536:25]
  assign outTag = ~inPipe_bits_singleOut; // @[FPU.scala 547:16]
  assign _T_54 = inPipe_bits_wflags & ~inPipe_bits_ren2; // @[FPU.scala 555:24]
  assign _T_57 = _T_8 ? 65'he008000000000000 : inPipe_bits_in1; // @[FPU.scala 558:24]
  assign fsgnjMux_data = _T_54 ? _T_57 : _GEN_23; // @[FPU.scala 555:42]
  assign _T_36 = {fsgnjMux_data[51:0], 24'h0}; // @[FPU.scala 231:28]
  assign _T_40 = fsgnjMux_data[63:52] + 12'h100; // @[FPU.scala 234:31]
  assign _T_42 = _T_40 - 12'h800; // @[FPU.scala 234:48]
  assign _T_43 = fsgnjMux_data[63:61] == 3'h0; // @[FPU.scala 235:19]
  assign _T_44 = fsgnjMux_data[63:61] >= 3'h6; // @[FPU.scala 235:36]
  assign _T_45 = _T_43 | _T_44; // @[FPU.scala 235:25]
  assign _T_47 = {fsgnjMux_data[63:61],_T_42[5:0]}; // @[Cat.scala 29:58]
  assign _T_49 = _T_45 ? _T_47 : _T_42[8:0]; // @[FPU.scala 235:10]
  assign _T_52 = {fsgnjMux_data[64:33],fsgnjMux_data[64],_T_49,_T_36[75:53]}; // @[Cat.scala 29:58]
  assign _T_63 = {_T_15, 4'h0}; // @[FPU.scala 560:51]
  assign _T_69 = {fsgnjMux_data[64:33],RecFNToRecFN_io_out}; // @[Cat.scala 29:58]
  assign io_out_bits_data = _T_71_data; // @[FPU.scala 577:10]
  assign io_out_bits_exc = _T_71_exc; // @[FPU.scala 577:10]
  assign RecFNToRecFN_io_in = inPipe_bits_in1; // @[FPU.scala 567:24]
  assign RecFNToRecFN_io_roundingMode = inPipe_bits_rm; // @[FPU.scala 568:34]
  assign FPToFP_cov_read_addr = FPToFP_state;
  assign FPToFP_cov_read_data = FPToFP_cov[FPToFP_cov_read_addr]; // @[Coverage map for FPToFP]
  assign FPToFP_cov_write_data = 1'h1;
  assign FPToFP_cov_write_addr = FPToFP_state;
  assign FPToFP_cov_write_mask = 1'h1;
  assign FPToFP_cov_write_en = 1'h1;
  assign inPipe_valid_shl = inPipe_valid;
  assign inPipe_valid_pad = {6'h0,inPipe_valid_shl};
  assign inPipe_bits_singleOut_shl = {inPipe_bits_singleOut, 1'h0};
  assign inPipe_bits_singleOut_pad = {5'h0,inPipe_bits_singleOut_shl};
  assign inPipe_bits_ren2_shl = {inPipe_bits_ren2, 2'h0};
  assign inPipe_bits_ren2_pad = {4'h0,inPipe_bits_ren2_shl};
  assign inPipe_bits_wflags_shl = {inPipe_bits_wflags, 3'h0};
  assign inPipe_bits_wflags_pad = {3'h0,inPipe_bits_wflags_shl};
  assign inPipe_bits_rm_shl = {inPipe_bits_rm, 4'h0};
  assign inPipe_bits_rm_pad = inPipe_bits_rm_shl;
  assign FPToFP_xor1 = inPipe_valid_pad ^ inPipe_bits_singleOut_pad;
  assign FPToFP_xor6 = inPipe_bits_wflags_pad ^ inPipe_bits_rm_pad;
  assign FPToFP_xor2 = inPipe_bits_ren2_pad ^ FPToFP_xor6;
  assign FPToFP_xor0 = FPToFP_xor1 ^ FPToFP_xor2;
  assign RecFNToRecFN_sum = FPToFP_covSum + RecFNToRecFN_io_covSum;
  assign io_covSum = RecFNToRecFN_sum;
  assign RecFNToRecFN_metaAssert_wire = RecFNToRecFN_metaAssert;
  assign metaAssert = FPToFP_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inPipe_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inPipe_bits_ren2 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  inPipe_bits_singleOut = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  inPipe_bits_wflags = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  inPipe_bits_rm = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  inPipe_bits_in1 = _RAND_5[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  inPipe_bits_in2 = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {3{`RANDOM}};
  _T_71_data = _RAND_7[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_71_exc = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  FPToFP_state = _RAND_9[6:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    FPToFP_cov[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  FPToFP_covSum = _RAND_11[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  FPToFP_metaAssert = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      inPipe_valid <= 1'h0;
    end else if (reset) begin
      inPipe_valid <= 1'h0;
    end else begin
      inPipe_valid <= io_in_valid;
    end
    if (metaReset) begin
      inPipe_bits_ren2 <= 1'h0;
    end else if (io_in_valid) begin
      inPipe_bits_ren2 <= io_in_bits_ren2;
    end
    if (metaReset) begin
      inPipe_bits_singleOut <= 1'h0;
    end else if (io_in_valid) begin
      inPipe_bits_singleOut <= io_in_bits_singleOut;
    end
    if (metaReset) begin
      inPipe_bits_wflags <= 1'h0;
    end else if (io_in_valid) begin
      inPipe_bits_wflags <= io_in_bits_wflags;
    end
    if (metaReset) begin
      inPipe_bits_rm <= 3'h0;
    end else if (io_in_valid) begin
      inPipe_bits_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      inPipe_bits_in1 <= 65'h0;
    end else if (io_in_valid) begin
      inPipe_bits_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      inPipe_bits_in2 <= 65'h0;
    end else if (io_in_valid) begin
      inPipe_bits_in2 <= io_in_bits_in2;
    end
    if (metaReset) begin
      _T_71_data <= 65'h0;
    end else if (inPipe_valid) begin
      if (_T_54) begin
        if (~outTag) begin
          _T_71_data <= _T_69;
        end else if (~outTag) begin
          _T_71_data <= _T_52;
        end else if (_T_54) begin
          if (_T_8) begin
            _T_71_data <= 65'he008000000000000;
          end else begin
            _T_71_data <= inPipe_bits_in1;
          end
        end else if (inPipe_bits_wflags) begin
          if (_T_22) begin
            _T_71_data <= 65'he008000000000000;
          end else if (_T_27) begin
            _T_71_data <= inPipe_bits_in1;
          end else begin
            _T_71_data <= inPipe_bits_in2;
          end
        end else begin
          _T_71_data <= fsgnj;
        end
      end else if (~outTag) begin
        _T_71_data <= _T_52;
      end else if (_T_54) begin
        if (_T_8) begin
          _T_71_data <= 65'he008000000000000;
        end else begin
          _T_71_data <= inPipe_bits_in1;
        end
      end else if (inPipe_bits_wflags) begin
        if (_T_22) begin
          _T_71_data <= 65'he008000000000000;
        end else if (_T_27) begin
          _T_71_data <= inPipe_bits_in1;
        end else begin
          _T_71_data <= inPipe_bits_in2;
        end
      end else begin
        _T_71_data <= fsgnj;
      end
    end
    if (metaReset) begin
      _T_71_exc <= 5'h0;
    end else if (inPipe_valid) begin
      if (_T_54) begin
        if (~outTag) begin
          _T_71_exc <= RecFNToRecFN_io_exceptionFlags;
        end else if (_T_54) begin
          _T_71_exc <= _T_63;
        end else if (inPipe_bits_wflags) begin
          _T_71_exc <= _T_28;
        end else begin
          _T_71_exc <= 5'h0;
        end
      end else if (_T_54) begin
        _T_71_exc <= _T_63;
      end else if (inPipe_bits_wflags) begin
        _T_71_exc <= _T_28;
      end else begin
        _T_71_exc <= 5'h0;
      end
    end
    FPToFP_state <= FPToFP_xor0;
    if (!(FPToFP_cov_read_data)) begin
      FPToFP_covSum <= FPToFP_covSum + 1'h1;
    end
    if (metaReset) begin
      FPToFP_metaAssert <= 1'h0;
    end else begin
      FPToFP_metaAssert <= FPToFP_metaAssert | RecFNToRecFN_metaAssert_wire;
    end
  end
  always @(posedge clock) begin
    if(FPToFP_cov_write_en & FPToFP_cov_write_mask) begin
      FPToFP_cov[FPToFP_cov_write_addr] <= FPToFP_cov_write_data; // @[Coverage map for FPToFP]
    end
  end
endmodule
module FPUFMAPipe_1(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_ren3,
  input         io_in_bits_swap23,
  input  [2:0]  io_in_bits_rm,
  input  [1:0]  io_in_bits_fmaCmd,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output [64:0] io_out_bits_data,
  output [4:0]  io_out_bits_exc,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         fma_halt
);
  wire  fma_clock; // @[FPU.scala 664:19]
  wire  fma_reset; // @[FPU.scala 664:19]
  wire  fma_io_validin; // @[FPU.scala 664:19]
  wire [1:0] fma_io_op; // @[FPU.scala 664:19]
  wire [64:0] fma_io_a; // @[FPU.scala 664:19]
  wire [64:0] fma_io_b; // @[FPU.scala 664:19]
  wire [64:0] fma_io_c; // @[FPU.scala 664:19]
  wire [2:0] fma_io_roundingMode; // @[FPU.scala 664:19]
  wire [64:0] fma_io_out; // @[FPU.scala 664:19]
  wire [4:0] fma_io_exceptionFlags; // @[FPU.scala 664:19]
  wire  fma_io_validout; // @[FPU.scala 664:19]
  wire [29:0] fma_io_covSum; // @[FPU.scala 664:19]
  wire  fma_metaAssert; // @[FPU.scala 664:19]
  wire  fma_metaReset; // @[FPU.scala 664:19]
  reg  valid; // @[FPU.scala 652:18]
  reg [31:0] _RAND_0;
  reg [2:0] in_rm; // @[FPU.scala 653:15]
  reg [31:0] _RAND_1;
  reg [1:0] in_fmaCmd; // @[FPU.scala 653:15]
  reg [31:0] _RAND_2;
  reg [64:0] in_in1; // @[FPU.scala 653:15]
  reg [95:0] _RAND_3;
  reg [64:0] in_in2; // @[FPU.scala 653:15]
  reg [95:0] _RAND_4;
  reg [64:0] in_in3; // @[FPU.scala 653:15]
  reg [95:0] _RAND_5;
  wire [64:0] _T_1; // @[FPU.scala 656:32]
  wire [64:0] _T_3; // @[FPU.scala 656:50]
  wire  _T_4; // @[FPU.scala 661:21]
  wire [64:0] _T_7; // @[FPU.scala 361:25]
  wire  _T_9; // @[FPU.scala 203:56]
  reg [64:0] _T_12_data; // @[Reg.scala 15:16]
  reg [95:0] _RAND_6;
  reg [4:0] _T_12_exc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  wire [4:0] res_exc; // @[FPU.scala 673:17 FPU.scala 675:11]
  wire [29:0] FPUFMAPipe_1_covSum;
  wire [29:0] fma_sum;
  wire  fma_metaAssert_wire;
  reg  FPUFMAPipe_1_metaAssert;
  reg [31:0] _RAND_8;
  MulAddRecFNPipe_1 fma ( // @[FPU.scala 664:19]
    .clock(fma_clock),
    .reset(fma_reset),
    .io_validin(fma_io_validin),
    .io_op(fma_io_op),
    .io_a(fma_io_a),
    .io_b(fma_io_b),
    .io_c(fma_io_c),
    .io_roundingMode(fma_io_roundingMode),
    .io_out(fma_io_out),
    .io_exceptionFlags(fma_io_exceptionFlags),
    .io_validout(fma_io_validout),
    .io_covSum(fma_io_covSum),
    .metaAssert(fma_metaAssert),
    .metaReset(fma_metaReset)
  );
  assign _T_1 = io_in_bits_in1 ^ io_in_bits_in2; // @[FPU.scala 656:32]
  assign _T_3 = _T_1 & 65'h10000000000000000; // @[FPU.scala 656:50]
  assign _T_4 = io_in_bits_ren3 | io_in_bits_swap23; // @[FPU.scala 661:21]
  assign _T_7 = fma_io_out & 65'h1efefffffffffffff; // @[FPU.scala 361:25]
  assign _T_9 = &fma_io_out[63:61]; // @[FPU.scala 203:56]
  assign res_exc = fma_io_exceptionFlags; // @[FPU.scala 673:17 FPU.scala 675:11]
  assign io_out_bits_data = _T_12_data; // @[FPU.scala 677:10]
  assign io_out_bits_exc = _T_12_exc; // @[FPU.scala 677:10]
  assign fma_clock = clock;
  assign fma_reset = reset;
  assign fma_io_validin = valid; // @[FPU.scala 665:18]
  assign fma_io_op = in_fmaCmd; // @[FPU.scala 666:13]
  assign fma_io_a = in_in1; // @[FPU.scala 669:12]
  assign fma_io_b = in_in2; // @[FPU.scala 670:12]
  assign fma_io_c = in_in3; // @[FPU.scala 671:12]
  assign fma_io_roundingMode = in_rm; // @[FPU.scala 667:23]
  assign FPUFMAPipe_1_covSum = 30'h0;
  assign fma_sum = FPUFMAPipe_1_covSum + fma_io_covSum;
  assign io_covSum = fma_sum;
  assign fma_metaAssert_wire = fma_metaAssert;
  assign metaAssert = FPUFMAPipe_1_metaAssert;
  assign fma_metaReset = metaReset | fma_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_rm = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_fmaCmd = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {3{`RANDOM}};
  in_in1 = _RAND_3[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {3{`RANDOM}};
  in_in2 = _RAND_4[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  in_in3 = _RAND_5[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  _T_12_data = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_12_exc = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  FPUFMAPipe_1_metaAssert = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      valid <= 1'h0;
    end else begin
      valid <= io_in_valid;
    end
    if (metaReset) begin
      in_rm <= 3'h0;
    end else if (io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      in_fmaCmd <= 2'h0;
    end else if (io_in_valid) begin
      in_fmaCmd <= io_in_bits_fmaCmd;
    end
    if (metaReset) begin
      in_in1 <= 65'h0;
    end else if (io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      in_in2 <= 65'h0;
    end else if (io_in_valid) begin
      if (io_in_bits_swap23) begin
        in_in2 <= 65'h8000000000000000;
      end else begin
        in_in2 <= io_in_bits_in2;
      end
    end
    if (metaReset) begin
      in_in3 <= 65'h0;
    end else if (io_in_valid) begin
      if (~_T_4) begin
        in_in3 <= _T_3;
      end else begin
        in_in3 <= io_in_bits_in3;
      end
    end
    if (metaReset) begin
      _T_12_data <= 65'h0;
    end else if (fma_io_validout) begin
      if (_T_9) begin
        _T_12_data <= _T_7;
      end else begin
        _T_12_data <= fma_io_out;
      end
    end
    if (metaReset) begin
      _T_12_exc <= 5'h0;
    end else if (fma_io_validout) begin
      _T_12_exc <= res_exc;
    end
    if (metaReset) begin
      FPUFMAPipe_1_metaAssert <= 1'h0;
    end else begin
      FPUFMAPipe_1_metaAssert <= FPUFMAPipe_1_metaAssert | fma_metaAssert_wire;
    end
  end
endmodule
module DivSqrtRecFN_small(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [2:0]  io_roundingMode,
  output        io_outValid_div,
  output        io_outValid_sqrt,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         divSqrtRecFNToRaw_halt
);
  wire  divSqrtRecFNToRaw_clock; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_reset; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_inValid; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_sqrtOp; // @[DivSqrtRecFN_small.scala 462:15]
  wire [32:0] divSqrtRecFNToRaw_io_a; // @[DivSqrtRecFN_small.scala 462:15]
  wire [32:0] divSqrtRecFNToRaw_io_b; // @[DivSqrtRecFN_small.scala 462:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingMode; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 462:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 462:15]
  wire [9:0] divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 462:15]
  wire [26:0] divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 462:15]
  wire [29:0] divSqrtRecFNToRaw_io_covSum; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_metaAssert; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_metaReset; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_divSqrtRawFN_halt; // @[DivSqrtRecFN_small.scala 462:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[DivSqrtRecFN_small.scala 477:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[DivSqrtRecFN_small.scala 477:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[DivSqrtRecFN_small.scala 477:15]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_detectTininess; // @[DivSqrtRecFN_small.scala 477:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 477:15]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 477:15]
  wire [29:0] roundRawFNToRecFN_io_covSum; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_metaAssert; // @[DivSqrtRecFN_small.scala 477:15]
  wire [29:0] DivSqrtRecFN_small_covSum;
  wire [29:0] divSqrtRecFNToRaw_sum;
  wire [29:0] roundRawFNToRecFN_sum;
  wire  divSqrtRecFNToRaw_metaAssert_wire;
  wire  roundRawFNToRecFN_metaAssert_wire;
  wire  DivSqrtRecFN_small_or0;
  reg  DivSqrtRecFN_small_metaAssert;
  reg [31:0] _RAND_0;
  DivSqrtRecFNToRaw_small divSqrtRecFNToRaw ( // @[DivSqrtRecFN_small.scala 462:15]
    .clock(divSqrtRecFNToRaw_clock),
    .reset(divSqrtRecFNToRaw_reset),
    .io_inReady(divSqrtRecFNToRaw_io_inReady),
    .io_inValid(divSqrtRecFNToRaw_io_inValid),
    .io_sqrtOp(divSqrtRecFNToRaw_io_sqrtOp),
    .io_a(divSqrtRecFNToRaw_io_a),
    .io_b(divSqrtRecFNToRaw_io_b),
    .io_roundingMode(divSqrtRecFNToRaw_io_roundingMode),
    .io_rawOutValid_div(divSqrtRecFNToRaw_io_rawOutValid_div),
    .io_rawOutValid_sqrt(divSqrtRecFNToRaw_io_rawOutValid_sqrt),
    .io_roundingModeOut(divSqrtRecFNToRaw_io_roundingModeOut),
    .io_invalidExc(divSqrtRecFNToRaw_io_invalidExc),
    .io_infiniteExc(divSqrtRecFNToRaw_io_infiniteExc),
    .io_rawOut_isNaN(divSqrtRecFNToRaw_io_rawOut_isNaN),
    .io_rawOut_isInf(divSqrtRecFNToRaw_io_rawOut_isInf),
    .io_rawOut_isZero(divSqrtRecFNToRaw_io_rawOut_isZero),
    .io_rawOut_sign(divSqrtRecFNToRaw_io_rawOut_sign),
    .io_rawOut_sExp(divSqrtRecFNToRaw_io_rawOut_sExp),
    .io_rawOut_sig(divSqrtRecFNToRaw_io_rawOut_sig),
    .io_covSum(divSqrtRecFNToRaw_io_covSum),
    .metaAssert(divSqrtRecFNToRaw_metaAssert),
    .metaReset(divSqrtRecFNToRaw_metaReset),
    .divSqrtRawFN_halt(divSqrtRecFNToRaw_divSqrtRawFN_halt)
  );
  RoundRawFNToRecFN_2 roundRawFNToRecFN ( // @[DivSqrtRecFN_small.scala 477:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundRawFNToRecFN_io_covSum),
    .metaAssert(roundRawFNToRecFN_metaAssert)
  );
  assign io_inReady = divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 464:16]
  assign io_outValid_div = divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 473:22]
  assign io_outValid_sqrt = divSqrtRecFNToRaw_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 474:22]
  assign io_out = roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 483:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 484:23]
  assign divSqrtRecFNToRaw_clock = clock;
  assign divSqrtRecFNToRaw_reset = reset;
  assign divSqrtRecFNToRaw_io_inValid = io_inValid; // @[DivSqrtRecFN_small.scala 465:39]
  assign divSqrtRecFNToRaw_io_sqrtOp = io_sqrtOp; // @[DivSqrtRecFN_small.scala 466:39]
  assign divSqrtRecFNToRaw_io_a = io_a; // @[DivSqrtRecFN_small.scala 467:39]
  assign divSqrtRecFNToRaw_io_b = io_b; // @[DivSqrtRecFN_small.scala 468:39]
  assign divSqrtRecFNToRaw_io_roundingMode = io_roundingMode; // @[DivSqrtRecFN_small.scala 469:39]
  assign roundRawFNToRecFN_io_invalidExc = divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 478:39]
  assign roundRawFNToRecFN_io_infiniteExc = divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 479:39]
  assign roundRawFNToRecFN_io_in_isNaN = divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_isInf = divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_isZero = divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_sign = divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_sExp = divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_sig = divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_roundingMode = divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 481:39]
  assign roundRawFNToRecFN_io_detectTininess = 1'h1; // @[DivSqrtRecFN_small.scala 482:41]
  assign DivSqrtRecFN_small_covSum = 30'h0;
  assign divSqrtRecFNToRaw_sum = DivSqrtRecFN_small_covSum + divSqrtRecFNToRaw_io_covSum;
  assign roundRawFNToRecFN_sum = divSqrtRecFNToRaw_sum + roundRawFNToRecFN_io_covSum;
  assign io_covSum = roundRawFNToRecFN_sum;
  assign divSqrtRecFNToRaw_metaAssert_wire = divSqrtRecFNToRaw_metaAssert;
  assign roundRawFNToRecFN_metaAssert_wire = roundRawFNToRecFN_metaAssert;
  assign DivSqrtRecFN_small_or0 = divSqrtRecFNToRaw_metaAssert_wire | roundRawFNToRecFN_metaAssert_wire;
  assign metaAssert = DivSqrtRecFN_small_metaAssert;
  assign divSqrtRecFNToRaw_metaReset = metaReset | divSqrtRecFNToRaw_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DivSqrtRecFN_small_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      DivSqrtRecFN_small_metaAssert <= 1'h0;
    end else begin
      DivSqrtRecFN_small_metaAssert <= DivSqrtRecFN_small_metaAssert | DivSqrtRecFN_small_or0;
    end
  end
endmodule
module DivSqrtRecFN_small_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [2:0]  io_roundingMode,
  output        io_outValid_div,
  output        io_outValid_sqrt,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         divSqrtRecFNToRaw_halt
);
  wire  divSqrtRecFNToRaw_clock; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_reset; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_inValid; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_sqrtOp; // @[DivSqrtRecFN_small.scala 462:15]
  wire [64:0] divSqrtRecFNToRaw_io_a; // @[DivSqrtRecFN_small.scala 462:15]
  wire [64:0] divSqrtRecFNToRaw_io_b; // @[DivSqrtRecFN_small.scala 462:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingMode; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 462:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 462:15]
  wire [12:0] divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 462:15]
  wire [55:0] divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 462:15]
  wire [29:0] divSqrtRecFNToRaw_io_covSum; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_metaAssert; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_metaReset; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_divSqrtRawFN_halt; // @[DivSqrtRecFN_small.scala 462:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[DivSqrtRecFN_small.scala 477:15]
  wire [12:0] roundRawFNToRecFN_io_in_sExp; // @[DivSqrtRecFN_small.scala 477:15]
  wire [55:0] roundRawFNToRecFN_io_in_sig; // @[DivSqrtRecFN_small.scala 477:15]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_detectTininess; // @[DivSqrtRecFN_small.scala 477:15]
  wire [64:0] roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 477:15]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 477:15]
  wire [29:0] roundRawFNToRecFN_io_covSum; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_metaAssert; // @[DivSqrtRecFN_small.scala 477:15]
  wire [29:0] DivSqrtRecFN_small_1_covSum;
  wire [29:0] divSqrtRecFNToRaw_sum;
  wire [29:0] roundRawFNToRecFN_sum;
  wire  divSqrtRecFNToRaw_metaAssert_wire;
  wire  roundRawFNToRecFN_metaAssert_wire;
  wire  DivSqrtRecFN_small_1_or0;
  reg  DivSqrtRecFN_small_1_metaAssert;
  reg [31:0] _RAND_0;
  DivSqrtRecFNToRaw_small_1 divSqrtRecFNToRaw ( // @[DivSqrtRecFN_small.scala 462:15]
    .clock(divSqrtRecFNToRaw_clock),
    .reset(divSqrtRecFNToRaw_reset),
    .io_inReady(divSqrtRecFNToRaw_io_inReady),
    .io_inValid(divSqrtRecFNToRaw_io_inValid),
    .io_sqrtOp(divSqrtRecFNToRaw_io_sqrtOp),
    .io_a(divSqrtRecFNToRaw_io_a),
    .io_b(divSqrtRecFNToRaw_io_b),
    .io_roundingMode(divSqrtRecFNToRaw_io_roundingMode),
    .io_rawOutValid_div(divSqrtRecFNToRaw_io_rawOutValid_div),
    .io_rawOutValid_sqrt(divSqrtRecFNToRaw_io_rawOutValid_sqrt),
    .io_roundingModeOut(divSqrtRecFNToRaw_io_roundingModeOut),
    .io_invalidExc(divSqrtRecFNToRaw_io_invalidExc),
    .io_infiniteExc(divSqrtRecFNToRaw_io_infiniteExc),
    .io_rawOut_isNaN(divSqrtRecFNToRaw_io_rawOut_isNaN),
    .io_rawOut_isInf(divSqrtRecFNToRaw_io_rawOut_isInf),
    .io_rawOut_isZero(divSqrtRecFNToRaw_io_rawOut_isZero),
    .io_rawOut_sign(divSqrtRecFNToRaw_io_rawOut_sign),
    .io_rawOut_sExp(divSqrtRecFNToRaw_io_rawOut_sExp),
    .io_rawOut_sig(divSqrtRecFNToRaw_io_rawOut_sig),
    .io_covSum(divSqrtRecFNToRaw_io_covSum),
    .metaAssert(divSqrtRecFNToRaw_metaAssert),
    .metaReset(divSqrtRecFNToRaw_metaReset),
    .divSqrtRawFN_halt(divSqrtRecFNToRaw_divSqrtRawFN_halt)
  );
  RoundRawFNToRecFN_3 roundRawFNToRecFN ( // @[DivSqrtRecFN_small.scala 477:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundRawFNToRecFN_io_covSum),
    .metaAssert(roundRawFNToRecFN_metaAssert)
  );
  assign io_inReady = divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 464:16]
  assign io_outValid_div = divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 473:22]
  assign io_outValid_sqrt = divSqrtRecFNToRaw_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 474:22]
  assign io_out = roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 483:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 484:23]
  assign divSqrtRecFNToRaw_clock = clock;
  assign divSqrtRecFNToRaw_reset = reset;
  assign divSqrtRecFNToRaw_io_inValid = io_inValid; // @[DivSqrtRecFN_small.scala 465:39]
  assign divSqrtRecFNToRaw_io_sqrtOp = io_sqrtOp; // @[DivSqrtRecFN_small.scala 466:39]
  assign divSqrtRecFNToRaw_io_a = io_a; // @[DivSqrtRecFN_small.scala 467:39]
  assign divSqrtRecFNToRaw_io_b = io_b; // @[DivSqrtRecFN_small.scala 468:39]
  assign divSqrtRecFNToRaw_io_roundingMode = io_roundingMode; // @[DivSqrtRecFN_small.scala 469:39]
  assign roundRawFNToRecFN_io_invalidExc = divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 478:39]
  assign roundRawFNToRecFN_io_infiniteExc = divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 479:39]
  assign roundRawFNToRecFN_io_in_isNaN = divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_isInf = divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_isZero = divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_sign = divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_sExp = divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_sig = divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_roundingMode = divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 481:39]
  assign roundRawFNToRecFN_io_detectTininess = 1'h1; // @[DivSqrtRecFN_small.scala 482:41]
  assign DivSqrtRecFN_small_1_covSum = 30'h0;
  assign divSqrtRecFNToRaw_sum = DivSqrtRecFN_small_1_covSum + divSqrtRecFNToRaw_io_covSum;
  assign roundRawFNToRecFN_sum = divSqrtRecFNToRaw_sum + roundRawFNToRecFN_io_covSum;
  assign io_covSum = roundRawFNToRecFN_sum;
  assign divSqrtRecFNToRaw_metaAssert_wire = divSqrtRecFNToRaw_metaAssert;
  assign roundRawFNToRecFN_metaAssert_wire = roundRawFNToRecFN_metaAssert;
  assign DivSqrtRecFN_small_1_or0 = divSqrtRecFNToRaw_metaAssert_wire | roundRawFNToRecFN_metaAssert_wire;
  assign metaAssert = DivSqrtRecFN_small_1_metaAssert;
  assign divSqrtRecFNToRaw_metaReset = metaReset | divSqrtRecFNToRaw_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DivSqrtRecFN_small_1_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      DivSqrtRecFN_small_1_metaAssert <= 1'h0;
    end else begin
      DivSqrtRecFN_small_1_metaAssert <= DivSqrtRecFN_small_1_metaAssert | DivSqrtRecFN_small_1_or0;
    end
  end
endmodule
module Arbiter(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [26:0] io_in_0_bits_bits_addr,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input         io_in_1_bits_valid,
  input  [26:0] io_in_1_bits_bits_addr,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_valid,
  output [26:0] io_out_bits_bits_addr,
  output        io_chosen,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  grant_1; // @[Arbiter.scala 31:78]
  wire [29:0] Arbiter_covSum;
  assign grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_valid = io_in_0_valid | io_in_1_bits_valid; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_bits_addr = io_in_0_valid ? io_in_0_bits_bits_addr : io_in_1_bits_bits_addr; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_chosen = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 123:13 Arbiter.scala 127:17]
  assign Arbiter_covSum = 30'h0;
  assign io_covSum = Arbiter_covSum;
  assign metaAssert = 1'h0;
endmodule
module OptimizationBarrier_117(
  input  [2:0]  io_x,
  output [2:0]  io_y,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] OptimizationBarrier_117_covSum;
  assign io_y = io_x; // @[package.scala 241:12]
  assign OptimizationBarrier_117_covSum = 30'h0;
  assign io_covSum = OptimizationBarrier_117_covSum;
  assign metaAssert = 1'h0;
endmodule
module OptimizationBarrier_118(
  input  [53:0] io_x_ppn,
  input         io_x_d,
  input         io_x_a,
  input         io_x_g,
  input         io_x_u,
  input         io_x_x,
  input         io_x_w,
  input         io_x_r,
  input         io_x_v,
  output [53:0] io_y_ppn,
  output        io_y_d,
  output        io_y_a,
  output        io_y_g,
  output        io_y_u,
  output        io_y_x,
  output        io_y_w,
  output        io_y_r,
  output        io_y_v,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] OptimizationBarrier_118_covSum;
  assign io_y_ppn = io_x_ppn; // @[package.scala 241:12]
  assign io_y_d = io_x_d; // @[package.scala 241:12]
  assign io_y_a = io_x_a; // @[package.scala 241:12]
  assign io_y_g = io_x_g; // @[package.scala 241:12]
  assign io_y_u = io_x_u; // @[package.scala 241:12]
  assign io_y_x = io_x_x; // @[package.scala 241:12]
  assign io_y_w = io_x_w; // @[package.scala 241:12]
  assign io_y_r = io_x_r; // @[package.scala 241:12]
  assign io_y_v = io_x_v; // @[package.scala 241:12]
  assign OptimizationBarrier_118_covSum = 30'h0;
  assign io_covSum = OptimizationBarrier_118_covSum;
  assign metaAssert = 1'h0;
endmodule
module IBuf(
  input         clock,
  input         reset,
  output        io_imem_ready,
  input         io_imem_valid,
  input         io_imem_bits_btb_taken,
  input         io_imem_bits_btb_bridx,
  input  [4:0]  io_imem_bits_btb_entry,
  input  [7:0]  io_imem_bits_btb_bht_history,
  input  [39:0] io_imem_bits_pc,
  input  [31:0] io_imem_bits_data,
  input         io_imem_bits_xcpt_pf_inst,
  input         io_imem_bits_xcpt_ae_inst,
  input         io_imem_bits_replay,
  input         io_kill,
  output [39:0] io_pc,
  output [4:0]  io_btb_resp_entry,
  output [7:0]  io_btb_resp_bht_history,
  input         io_inst_0_ready,
  output        io_inst_0_valid,
  output        io_inst_0_bits_xcpt0_pf_inst,
  output        io_inst_0_bits_xcpt0_ae_inst,
  output        io_inst_0_bits_xcpt1_pf_inst,
  output        io_inst_0_bits_xcpt1_ae_inst,
  output        io_inst_0_bits_replay,
  output        io_inst_0_bits_rvc,
  output [31:0] io_inst_0_bits_inst_bits,
  output [4:0]  io_inst_0_bits_inst_rd,
  output [4:0]  io_inst_0_bits_inst_rs1,
  output [4:0]  io_inst_0_bits_inst_rs2,
  output [4:0]  io_inst_0_bits_inst_rs3,
  output [31:0] io_inst_0_bits_raw,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [31:0] RVCExpander_io_in; // @[IBuf.scala 86:21]
  wire [31:0] RVCExpander_io_out_bits; // @[IBuf.scala 86:21]
  wire [4:0] RVCExpander_io_out_rd; // @[IBuf.scala 86:21]
  wire [4:0] RVCExpander_io_out_rs1; // @[IBuf.scala 86:21]
  wire [4:0] RVCExpander_io_out_rs2; // @[IBuf.scala 86:21]
  wire [4:0] RVCExpander_io_out_rs3; // @[IBuf.scala 86:21]
  wire  RVCExpander_io_rvc; // @[IBuf.scala 86:21]
  wire [29:0] RVCExpander_io_covSum; // @[IBuf.scala 86:21]
  wire  RVCExpander_metaAssert; // @[IBuf.scala 86:21]
  reg  nBufValid; // @[IBuf.scala 34:47]
  reg [31:0] _RAND_0;
  reg [39:0] buf__pc; // @[IBuf.scala 35:16]
  reg [63:0] _RAND_1;
  reg [31:0] buf__data; // @[IBuf.scala 35:16]
  reg [31:0] _RAND_2;
  reg  buf__xcpt_pf_inst; // @[IBuf.scala 35:16]
  reg [31:0] _RAND_3;
  reg  buf__xcpt_ae_inst; // @[IBuf.scala 35:16]
  reg [31:0] _RAND_4;
  reg  buf__replay; // @[IBuf.scala 35:16]
  reg [31:0] _RAND_5;
  reg [4:0] ibufBTBResp_entry; // @[IBuf.scala 36:24]
  reg [31:0] _RAND_6;
  reg [7:0] ibufBTBResp_bht_history; // @[IBuf.scala 36:24]
  reg [31:0] _RAND_7;
  wire  pcWordBits; // @[package.scala 143:13]
  wire [1:0] _T; // @[IBuf.scala 41:64]
  wire [1:0] _T_1; // @[IBuf.scala 41:16]
  wire [1:0] _GEN_56; // @[IBuf.scala 41:88]
  wire [1:0] nIC; // @[IBuf.scala 41:88]
  wire [1:0] _T_4; // @[IBuf.scala 43:19]
  wire [1:0] _GEN_57; // @[IBuf.scala 43:49]
  wire [1:0] nValid; // @[IBuf.scala 43:49]
  wire [3:0] _T_62; // @[OneHot.scala 58:35]
  wire [3:0] _T_64; // @[IBuf.scala 74:33]
  wire [1:0] valid; // @[IBuf.scala 74:37]
  wire [1:0] _T_93; // @[IBuf.scala 93:42]
  wire  _T_95; // @[IBuf.scala 93:34]
  wire [1:0] _T_65; // @[OneHot.scala 58:35]
  wire [1:0] bufMask; // @[IBuf.scala 75:37]
  wire [1:0] buf_replay; // @[IBuf.scala 77:23]
  wire  _T_98; // @[IBuf.scala 93:48]
  wire [1:0] _T_128; // @[IBuf.scala 102:71]
  wire [1:0] nReady; // @[IBuf.scala 102:56]
  wire [1:0] nICReady; // @[IBuf.scala 42:25]
  wire  _T_6; // @[IBuf.scala 44:47]
  wire  _T_7; // @[IBuf.scala 44:37]
  wire  _T_8; // @[IBuf.scala 44:73]
  wire [1:0] _T_10; // @[IBuf.scala 44:92]
  wire  _T_11; // @[IBuf.scala 44:85]
  wire  _T_12; // @[IBuf.scala 44:80]
  wire [1:0] _T_16; // @[IBuf.scala 48:64]
  wire [1:0] _T_17; // @[IBuf.scala 48:23]
  wire  _T_19; // @[IBuf.scala 54:27]
  wire  _T_20; // @[IBuf.scala 54:62]
  wire  _T_21; // @[IBuf.scala 54:50]
  wire  _T_25; // @[IBuf.scala 54:68]
  wire [1:0] _T_27; // @[IBuf.scala 55:32]
  wire [63:0] _T_32; // @[Cat.scala 29:58]
  wire [5:0] _T_33; // @[IBuf.scala 128:19]
  wire [63:0] _T_34; // @[IBuf.scala 128:10]
  wire [39:0] _T_37; // @[IBuf.scala 59:35]
  wire [2:0] _T_38; // @[IBuf.scala 59:80]
  wire [39:0] _GEN_65; // @[IBuf.scala 59:68]
  wire [39:0] _T_40; // @[IBuf.scala 59:68]
  wire [39:0] _T_41; // @[IBuf.scala 59:109]
  wire [39:0] _T_42; // @[IBuf.scala 59:49]
  wire [1:0] _GEN_0; // @[IBuf.scala 54:92]
  wire [1:0] _GEN_23; // @[IBuf.scala 47:29]
  wire [1:0] _GEN_46; // @[IBuf.scala 63:20]
  wire [1:0] _T_44; // @[IBuf.scala 68:32]
  wire [1:0] icShiftAmt; // @[IBuf.scala 68:44]
  wire [63:0] _T_49; // @[Cat.scala 29:58]
  wire [127:0] _T_53; // @[Cat.scala 29:58]
  wire [5:0] _T_54; // @[IBuf.scala 121:19]
  wire [190:0] _GEN_68; // @[IBuf.scala 121:10]
  wire [190:0] _T_55; // @[IBuf.scala 121:10]
  wire [31:0] icData; // @[package.scala 143:13]
  wire [4:0] _T_57; // @[IBuf.scala 71:65]
  wire [62:0] _T_58; // @[IBuf.scala 71:51]
  wire [31:0] icMask; // @[IBuf.scala 71:92]
  wire [31:0] _T_59; // @[IBuf.scala 72:21]
  wire [31:0] _T_61; // @[IBuf.scala 72:41]
  wire  xcpt_1_pf_inst; // @[IBuf.scala 76:53]
  wire  xcpt_1_ae_inst; // @[IBuf.scala 76:53]
  wire [1:0] _T_70; // @[IBuf.scala 78:63]
  wire [1:0] _T_71; // @[IBuf.scala 78:35]
  wire [1:0] ic_replay; // @[IBuf.scala 78:30]
  wire  _T_74; // @[IBuf.scala 79:25]
  wire  _T_75; // @[IBuf.scala 79:78]
  wire  _T_76; // @[IBuf.scala 79:52]
  wire  _T_78; // @[IBuf.scala 79:9]
  wire  _T_80; // @[IBuf.scala 82:26]
  wire [1:0] _T_87; // @[IBuf.scala 92:61]
  wire  _T_89; // @[IBuf.scala 92:49]
  wire [1:0] _T_108; // @[IBuf.scala 96:63]
  wire [1:0] _T_109; // @[IBuf.scala 96:35]
  wire  _T_116; // @[IBuf.scala 100:25]
  wire [1:0] _T_119; // @[IBuf.scala 100:50]
  wire  _T_121; // @[IBuf.scala 100:40]
  reg [1:0] IBuf_state; // @[Register tracking IBuf state]
  reg [31:0] _RAND_8;
  reg  IBuf_cov [0:3]; // @[Coverage map for IBuf]
  reg [31:0] _RAND_9;
  wire  IBuf_cov_read_data; // @[Coverage map for IBuf]
  wire [1:0] IBuf_cov_read_addr; // @[Coverage map for IBuf]
  wire  IBuf_cov_write_data; // @[Coverage map for IBuf]
  wire [1:0] IBuf_cov_write_addr; // @[Coverage map for IBuf]
  wire  IBuf_cov_write_mask; // @[Coverage map for IBuf]
  wire  IBuf_cov_write_en; // @[Coverage map for IBuf]
  reg [29:0] IBuf_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_10;
  wire  nBufValid_shl;
  wire [1:0] nBufValid_pad;
  wire [1:0] buf__replay_shl;
  wire [1:0] buf__replay_pad;
  wire [1:0] IBuf_xor0;
  wire [29:0] RVCExpander_sum;
  wire  stopEn0;
  wire  RVCExpander_metaAssert_wire;
  wire  IBuf_or0;
  reg  IBuf_metaAssert;
  reg [31:0] _RAND_11;
  RVCExpander RVCExpander ( // @[IBuf.scala 86:21]
    .io_in(RVCExpander_io_in),
    .io_out_bits(RVCExpander_io_out_bits),
    .io_out_rd(RVCExpander_io_out_rd),
    .io_out_rs1(RVCExpander_io_out_rs1),
    .io_out_rs2(RVCExpander_io_out_rs2),
    .io_out_rs3(RVCExpander_io_out_rs3),
    .io_rvc(RVCExpander_io_rvc),
    .io_covSum(RVCExpander_io_covSum),
    .metaAssert(RVCExpander_metaAssert)
  );
  assign pcWordBits = io_imem_bits_pc[1]; // @[package.scala 143:13]
  assign _T = io_imem_bits_btb_bridx + 1'h1; // @[IBuf.scala 41:64]
  assign _T_1 = io_imem_bits_btb_taken ? _T : 2'h2; // @[IBuf.scala 41:16]
  assign _GEN_56 = {{1'd0}, pcWordBits}; // @[IBuf.scala 41:88]
  assign nIC = _T_1 - _GEN_56; // @[IBuf.scala 41:88]
  assign _T_4 = io_imem_valid ? nIC : 2'h0; // @[IBuf.scala 43:19]
  assign _GEN_57 = {{1'd0}, nBufValid}; // @[IBuf.scala 43:49]
  assign nValid = _T_4 + _GEN_57; // @[IBuf.scala 43:49]
  assign _T_62 = 4'h1 << nValid; // @[OneHot.scala 58:35]
  assign _T_64 = _T_62 - 4'h1; // @[IBuf.scala 74:33]
  assign valid = _T_64[1:0]; // @[IBuf.scala 74:37]
  assign _T_93 = {{1'd0}, valid[1]}; // @[IBuf.scala 93:42]
  assign _T_95 = RVCExpander_io_rvc | _T_93[0]; // @[IBuf.scala 93:34]
  assign _T_65 = 2'h1 << nBufValid; // @[OneHot.scala 58:35]
  assign bufMask = _T_65 - 2'h1; // @[IBuf.scala 75:37]
  assign buf_replay = buf__replay ? bufMask : 2'h0; // @[IBuf.scala 77:23]
  assign _T_98 = _T_95 | buf_replay[0]; // @[IBuf.scala 93:48]
  assign _T_128 = RVCExpander_io_rvc ? 2'h1 : 2'h2; // @[IBuf.scala 102:71]
  assign nReady = _T_98 ? _T_128 : 2'h0; // @[IBuf.scala 102:56]
  assign nICReady = nReady - _GEN_57; // @[IBuf.scala 42:25]
  assign _T_6 = nReady >= _GEN_57; // @[IBuf.scala 44:47]
  assign _T_7 = io_inst_0_ready & _T_6; // @[IBuf.scala 44:37]
  assign _T_8 = nICReady >= nIC; // @[IBuf.scala 44:73]
  assign _T_10 = nIC - nICReady; // @[IBuf.scala 44:92]
  assign _T_11 = 2'h1 >= _T_10; // @[IBuf.scala 44:85]
  assign _T_12 = _T_8 | _T_11; // @[IBuf.scala 44:80]
  assign _T_16 = _GEN_57 - nReady; // @[IBuf.scala 48:64]
  assign _T_17 = _T_6 ? 2'h0 : _T_16; // @[IBuf.scala 48:23]
  assign _T_19 = io_imem_valid & _T_6; // @[IBuf.scala 54:27]
  assign _T_20 = nICReady < nIC; // @[IBuf.scala 54:62]
  assign _T_21 = _T_19 & _T_20; // @[IBuf.scala 54:50]
  assign _T_25 = _T_21 & _T_11; // @[IBuf.scala 54:68]
  assign _T_27 = _GEN_56 + nICReady; // @[IBuf.scala 55:32]
  assign _T_32 = {io_imem_bits_data[31:16],io_imem_bits_data[31:16],io_imem_bits_data}; // @[Cat.scala 29:58]
  assign _T_33 = {_T_27, 4'h0}; // @[IBuf.scala 128:19]
  assign _T_34 = _T_32 >> _T_33; // @[IBuf.scala 128:10]
  assign _T_37 = io_imem_bits_pc & 40'hfffffffffc; // @[IBuf.scala 59:35]
  assign _T_38 = {nICReady, 1'h0}; // @[IBuf.scala 59:80]
  assign _GEN_65 = {{37'd0}, _T_38}; // @[IBuf.scala 59:68]
  assign _T_40 = io_imem_bits_pc + _GEN_65; // @[IBuf.scala 59:68]
  assign _T_41 = _T_40 & 40'h3; // @[IBuf.scala 59:109]
  assign _T_42 = _T_37 | _T_41; // @[IBuf.scala 59:49]
  assign _GEN_0 = _T_25 ? _T_10 : _T_17; // @[IBuf.scala 54:92]
  assign _GEN_23 = io_inst_0_ready ? _GEN_0 : {{1'd0}, nBufValid}; // @[IBuf.scala 47:29]
  assign _GEN_46 = io_kill ? 2'h0 : _GEN_23; // @[IBuf.scala 63:20]
  assign _T_44 = 2'h2 + _GEN_57; // @[IBuf.scala 68:32]
  assign icShiftAmt = _T_44 - _GEN_56; // @[IBuf.scala 68:44]
  assign _T_49 = {io_imem_bits_data,io_imem_bits_data[15:0],io_imem_bits_data[15:0]}; // @[Cat.scala 29:58]
  assign _T_53 = {_T_49[63:48],_T_49[63:48],_T_49[63:48],_T_49[63:48],io_imem_bits_data,io_imem_bits_data[15:0],io_imem_bits_data[15:0]}; // @[Cat.scala 29:58]
  assign _T_54 = {icShiftAmt, 4'h0}; // @[IBuf.scala 121:19]
  assign _GEN_68 = {{63'd0}, _T_53}; // @[IBuf.scala 121:10]
  assign _T_55 = _GEN_68 << _T_54; // @[IBuf.scala 121:10]
  assign icData = _T_55[95:64]; // @[package.scala 143:13]
  assign _T_57 = {nBufValid, 4'h0}; // @[IBuf.scala 71:65]
  assign _T_58 = 63'hffffffff << _T_57; // @[IBuf.scala 71:51]
  assign icMask = _T_58[31:0]; // @[IBuf.scala 71:92]
  assign _T_59 = icData & icMask; // @[IBuf.scala 72:21]
  assign _T_61 = buf__data & ~icMask; // @[IBuf.scala 72:41]
  assign xcpt_1_pf_inst = bufMask[1] ? buf__xcpt_pf_inst : io_imem_bits_xcpt_pf_inst; // @[IBuf.scala 76:53]
  assign xcpt_1_ae_inst = bufMask[1] ? buf__xcpt_ae_inst : io_imem_bits_xcpt_ae_inst; // @[IBuf.scala 76:53]
  assign _T_70 = valid & ~bufMask; // @[IBuf.scala 78:63]
  assign _T_71 = io_imem_bits_replay ? _T_70 : 2'h0; // @[IBuf.scala 78:35]
  assign ic_replay = buf_replay | _T_71; // @[IBuf.scala 78:30]
  assign _T_74 = ~io_imem_valid | ~io_imem_bits_btb_taken; // @[IBuf.scala 79:25]
  assign _T_75 = io_imem_bits_btb_bridx >= pcWordBits; // @[IBuf.scala 79:78]
  assign _T_76 = _T_74 | _T_75; // @[IBuf.scala 79:52]
  assign _T_78 = _T_76 | reset; // @[IBuf.scala 79:9]
  assign _T_80 = nBufValid > 1'h0; // @[IBuf.scala 82:26]
  assign _T_87 = {{1'd0}, ic_replay[1]}; // @[IBuf.scala 92:61]
  assign _T_89 = ~RVCExpander_io_rvc & _T_87[0]; // @[IBuf.scala 92:49]
  assign _T_108 = {xcpt_1_pf_inst,xcpt_1_ae_inst}; // @[IBuf.scala 96:63]
  assign _T_109 = RVCExpander_io_rvc ? 2'h0 : _T_108; // @[IBuf.scala 96:35]
  assign _T_116 = bufMask[0] & RVCExpander_io_rvc; // @[IBuf.scala 100:25]
  assign _T_119 = {{1'd0}, bufMask[1]}; // @[IBuf.scala 100:50]
  assign _T_121 = _T_116 | _T_119[0]; // @[IBuf.scala 100:40]
  assign io_imem_ready = _T_7 & _T_12; // @[IBuf.scala 44:17]
  assign io_pc = _T_80 ? buf__pc : io_imem_bits_pc; // @[IBuf.scala 82:9]
  assign io_btb_resp_entry = _T_121 ? ibufBTBResp_entry : io_imem_bits_btb_entry; // @[IBuf.scala 81:15 IBuf.scala 100:71]
  assign io_btb_resp_bht_history = _T_121 ? ibufBTBResp_bht_history : io_imem_bits_btb_bht_history; // @[IBuf.scala 81:15 IBuf.scala 100:71]
  assign io_inst_0_valid = valid[0] & _T_98; // @[IBuf.scala 94:24]
  assign io_inst_0_bits_xcpt0_pf_inst = bufMask[0] ? buf__xcpt_pf_inst : io_imem_bits_xcpt_pf_inst; // @[IBuf.scala 95:29]
  assign io_inst_0_bits_xcpt0_ae_inst = bufMask[0] ? buf__xcpt_ae_inst : io_imem_bits_xcpt_ae_inst; // @[IBuf.scala 95:29]
  assign io_inst_0_bits_xcpt1_pf_inst = _T_109[1]; // @[IBuf.scala 96:29]
  assign io_inst_0_bits_xcpt1_ae_inst = _T_109[0]; // @[IBuf.scala 96:29]
  assign io_inst_0_bits_replay = ic_replay[0] | _T_89; // @[IBuf.scala 97:30]
  assign io_inst_0_bits_rvc = RVCExpander_io_rvc; // @[IBuf.scala 98:27]
  assign io_inst_0_bits_inst_bits = RVCExpander_io_out_bits; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rd = RVCExpander_io_out_rd; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rs1 = RVCExpander_io_out_rs1; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rs2 = RVCExpander_io_out_rs2; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rs3 = RVCExpander_io_out_rs3; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_raw = _T_59 | _T_61; // @[IBuf.scala 89:25]
  assign RVCExpander_io_in = _T_59 | _T_61; // @[IBuf.scala 87:15]
  assign IBuf_cov_read_addr = IBuf_state;
  assign IBuf_cov_read_data = IBuf_cov[IBuf_cov_read_addr]; // @[Coverage map for IBuf]
  assign IBuf_cov_write_data = 1'h1;
  assign IBuf_cov_write_addr = IBuf_state;
  assign IBuf_cov_write_mask = 1'h1;
  assign IBuf_cov_write_en = 1'h1;
  assign nBufValid_shl = nBufValid;
  assign nBufValid_pad = {1'h0,nBufValid_shl};
  assign buf__replay_shl = {buf__replay, 1'h0};
  assign buf__replay_pad = buf__replay_shl;
  assign IBuf_xor0 = nBufValid_pad ^ buf__replay_pad;
  assign RVCExpander_sum = IBuf_covSum + RVCExpander_io_covSum;
  assign io_covSum = RVCExpander_sum;
  assign stopEn0 = ~_T_78;
  assign RVCExpander_metaAssert_wire = RVCExpander_metaAssert;
  assign IBuf_or0 = stopEn0 | RVCExpander_metaAssert_wire;
  assign metaAssert = IBuf_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  nBufValid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  buf__pc = _RAND_1[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  buf__data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  buf__xcpt_pf_inst = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  buf__xcpt_ae_inst = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  buf__replay = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ibufBTBResp_entry = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ibufBTBResp_bht_history = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  IBuf_state = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    IBuf_cov[initvar] = _RAND_9[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  IBuf_covSum = _RAND_10[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  IBuf_metaAssert = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      nBufValid <= 1'h0;
    end else if (reset) begin
      nBufValid <= 1'h0;
    end else begin
      nBufValid <= _GEN_46[0];
    end
    if (metaReset) begin
      buf__pc <= 40'h0;
    end else if (io_inst_0_ready) begin
      if (_T_25) begin
        buf__pc <= _T_42;
      end
    end
    if (metaReset) begin
      buf__data <= 32'h0;
    end else if (io_inst_0_ready) begin
      if (_T_25) begin
        buf__data <= {{16'd0}, _T_34[15:0]};
      end
    end
    if (metaReset) begin
      buf__xcpt_pf_inst <= 1'h0;
    end else if (io_inst_0_ready) begin
      if (_T_25) begin
        buf__xcpt_pf_inst <= io_imem_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      buf__xcpt_ae_inst <= 1'h0;
    end else if (io_inst_0_ready) begin
      if (_T_25) begin
        buf__xcpt_ae_inst <= io_imem_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      buf__replay <= 1'h0;
    end else if (io_inst_0_ready) begin
      if (_T_25) begin
        buf__replay <= io_imem_bits_replay;
      end
    end
    if (metaReset) begin
      ibufBTBResp_entry <= 5'h0;
    end else if (io_inst_0_ready) begin
      if (_T_25) begin
        ibufBTBResp_entry <= io_imem_bits_btb_entry;
      end
    end
    if (metaReset) begin
      ibufBTBResp_bht_history <= 8'h0;
    end else if (io_inst_0_ready) begin
      if (_T_25) begin
        ibufBTBResp_bht_history <= io_imem_bits_btb_bht_history;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_78) begin
          $fwrite(32'h80000002,"Assertion failed\n    at IBuf.scala:79 assert(!io.imem.valid || !io.imem.bits.btb.taken || io.imem.bits.btb.bridx >= pcWordBits)\n"); // @[IBuf.scala 79:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_78) begin
          $fatal; // @[IBuf.scala 79:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    IBuf_state <= IBuf_xor0;
    if (!(IBuf_cov_read_data)) begin
      IBuf_covSum <= IBuf_covSum + 1'h1;
    end
    if (metaReset) begin
      IBuf_metaAssert <= 1'h0;
    end else begin
      IBuf_metaAssert <= IBuf_metaAssert | IBuf_or0;
    end
  end
  always @(posedge clock) begin
    if(IBuf_cov_write_en & IBuf_cov_write_mask) begin
      IBuf_cov[IBuf_cov_write_addr] <= IBuf_cov_write_data; // @[Coverage map for IBuf]
    end
  end
endmodule
module CSRFile(
  input         clock,
  input         reset,
  input         io_ungated_clock,
  input         io_interrupts_debug,
  input         io_interrupts_mtip,
  input         io_interrupts_msip,
  input         io_interrupts_meip,
  input         io_interrupts_seip,
  input         io_hartid,
  input  [11:0] io_rw_addr,
  input  [2:0]  io_rw_cmd,
  output [63:0] io_rw_rdata,
  input  [63:0] io_rw_wdata,
  input  [11:0] io_decode_0_csr,
  output        io_decode_0_fp_illegal,
  output        io_decode_0_fp_csr,
  output        io_decode_0_read_illegal,
  output        io_decode_0_write_illegal,
  output        io_decode_0_write_flush,
  output        io_decode_0_system_illegal,
  output        io_csr_stall,
  output        io_eret,
  output        io_singleStep,
  output        io_status_debug,
  output        io_status_cease,
  output        io_status_wfi,
  output [31:0] io_status_isa,
  output [1:0]  io_status_dprv,
  output [1:0]  io_status_prv,
  output        io_status_sd,
  output [26:0] io_status_zero2,
  output [1:0]  io_status_sxl,
  output [1:0]  io_status_uxl,
  output        io_status_sd_rv32,
  output [7:0]  io_status_zero1,
  output        io_status_tsr,
  output        io_status_tw,
  output        io_status_tvm,
  output        io_status_mxr,
  output        io_status_sum,
  output        io_status_mprv,
  output [1:0]  io_status_xs,
  output [1:0]  io_status_fs,
  output [1:0]  io_status_mpp,
  output [1:0]  io_status_vs,
  output        io_status_spp,
  output        io_status_mpie,
  output        io_status_hpie,
  output        io_status_spie,
  output        io_status_upie,
  output        io_status_mie,
  output        io_status_hie,
  output        io_status_sie,
  output        io_status_uie,
  output [3:0]  io_ptbr_mode,
  output [43:0] io_ptbr_ppn,
  output [39:0] io_evec,
  input         io_exception,
  input         io_retire,
  input  [63:0] io_cause,
  input  [39:0] io_pc,
  input  [39:0] io_tval,
  output [63:0] io_time,
  output [2:0]  io_fcsr_rm,
  input         io_fcsr_flags_valid,
  input  [4:0]  io_fcsr_flags_bits,
  output        io_interrupt,
  output [63:0] io_interrupt_cause,
  output        io_bp_0_control_action,
  output [1:0]  io_bp_0_control_tmatch,
  output        io_bp_0_control_m,
  output        io_bp_0_control_s,
  output        io_bp_0_control_u,
  output        io_bp_0_control_x,
  output        io_bp_0_control_w,
  output        io_bp_0_control_r,
  output [38:0] io_bp_0_address,
  output        io_pmp_0_cfg_l,
  output [1:0]  io_pmp_0_cfg_a,
  output        io_pmp_0_cfg_x,
  output        io_pmp_0_cfg_w,
  output        io_pmp_0_cfg_r,
  output [29:0] io_pmp_0_addr,
  output [31:0] io_pmp_0_mask,
  output        io_pmp_1_cfg_l,
  output [1:0]  io_pmp_1_cfg_a,
  output        io_pmp_1_cfg_x,
  output        io_pmp_1_cfg_w,
  output        io_pmp_1_cfg_r,
  output [29:0] io_pmp_1_addr,
  output [31:0] io_pmp_1_mask,
  output        io_pmp_2_cfg_l,
  output [1:0]  io_pmp_2_cfg_a,
  output        io_pmp_2_cfg_x,
  output        io_pmp_2_cfg_w,
  output        io_pmp_2_cfg_r,
  output [29:0] io_pmp_2_addr,
  output [31:0] io_pmp_2_mask,
  output        io_pmp_3_cfg_l,
  output [1:0]  io_pmp_3_cfg_a,
  output        io_pmp_3_cfg_x,
  output        io_pmp_3_cfg_w,
  output        io_pmp_3_cfg_r,
  output [29:0] io_pmp_3_addr,
  output [31:0] io_pmp_3_mask,
  output        io_pmp_4_cfg_l,
  output [1:0]  io_pmp_4_cfg_a,
  output        io_pmp_4_cfg_x,
  output        io_pmp_4_cfg_w,
  output        io_pmp_4_cfg_r,
  output [29:0] io_pmp_4_addr,
  output [31:0] io_pmp_4_mask,
  output        io_pmp_5_cfg_l,
  output [1:0]  io_pmp_5_cfg_a,
  output        io_pmp_5_cfg_x,
  output        io_pmp_5_cfg_w,
  output        io_pmp_5_cfg_r,
  output [29:0] io_pmp_5_addr,
  output [31:0] io_pmp_5_mask,
  output        io_pmp_6_cfg_l,
  output [1:0]  io_pmp_6_cfg_a,
  output        io_pmp_6_cfg_x,
  output        io_pmp_6_cfg_w,
  output        io_pmp_6_cfg_r,
  output [29:0] io_pmp_6_addr,
  output [31:0] io_pmp_6_mask,
  output        io_pmp_7_cfg_l,
  output [1:0]  io_pmp_7_cfg_a,
  output        io_pmp_7_cfg_x,
  output        io_pmp_7_cfg_w,
  output        io_pmp_7_cfg_r,
  output [29:0] io_pmp_7_addr,
  output [31:0] io_pmp_7_mask,
  input  [31:0] io_inst_0,
  output        io_trace_0_valid,
  output [39:0] io_trace_0_iaddr,
  output [31:0] io_trace_0_insn,
  output        io_trace_0_exception,
  output [63:0] io_customCSRs_0_value,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [1:0] reg_mstatus_prv; // @[CSR.scala 312:24]
  reg [31:0] _RAND_0;
  reg  reg_mstatus_tsr; // @[CSR.scala 312:24]
  reg [31:0] _RAND_1;
  reg  reg_mstatus_tw; // @[CSR.scala 312:24]
  reg [31:0] _RAND_2;
  reg  reg_mstatus_tvm; // @[CSR.scala 312:24]
  reg [31:0] _RAND_3;
  reg  reg_mstatus_mxr; // @[CSR.scala 312:24]
  reg [31:0] _RAND_4;
  reg  reg_mstatus_sum; // @[CSR.scala 312:24]
  reg [31:0] _RAND_5;
  reg  reg_mstatus_mprv; // @[CSR.scala 312:24]
  reg [31:0] _RAND_6;
  reg [1:0] reg_mstatus_fs; // @[CSR.scala 312:24]
  reg [31:0] _RAND_7;
  reg [1:0] reg_mstatus_mpp; // @[CSR.scala 312:24]
  reg [31:0] _RAND_8;
  reg  reg_mstatus_spp; // @[CSR.scala 312:24]
  reg [31:0] _RAND_9;
  reg  reg_mstatus_mpie; // @[CSR.scala 312:24]
  reg [31:0] _RAND_10;
  reg  reg_mstatus_spie; // @[CSR.scala 312:24]
  reg [31:0] _RAND_11;
  reg  reg_mstatus_mie; // @[CSR.scala 312:24]
  reg [31:0] _RAND_12;
  reg  reg_mstatus_sie; // @[CSR.scala 312:24]
  reg [31:0] _RAND_13;
  wire  system_insn; // @[CSR.scala 589:31]
  wire [31:0] _T_703; // @[CSR.scala 601:28]
  wire [31:0] _T_710; // @[Decode.scala 14:65]
  wire  _T_711; // @[Decode.scala 14:121]
  wire [31:0] _T_712; // @[Decode.scala 14:65]
  wire  _T_713; // @[Decode.scala 14:121]
  wire  _T_715; // @[Decode.scala 15:30]
  wire  insn_ret; // @[CSR.scala 601:95]
  reg [1:0] reg_dcsr_prv; // @[CSR.scala 320:21]
  reg [31:0] _RAND_14;
  wire [1:0] _GEN_93; // @[CSR.scala 745:53]
  wire [1:0] _GEN_102; // @[CSR.scala 739:52]
  wire [31:0] _T_704; // @[Decode.scala 14:65]
  wire  _T_705; // @[Decode.scala 14:121]
  wire  insn_call; // @[CSR.scala 601:95]
  wire  _T_708; // @[Decode.scala 14:121]
  wire  insn_break; // @[CSR.scala 601:95]
  wire  _T_1197; // @[CSR.scala 673:29]
  wire  exception; // @[CSR.scala 673:43]
  reg  reg_singleStepped; // @[CSR.scala 364:30]
  reg [31:0] _RAND_15;
  wire [3:0] _GEN_490; // @[CSR.scala 637:36]
  wire [3:0] _T_1143; // @[CSR.scala 637:36]
  wire [63:0] _T_1144; // @[CSR.scala 638:14]
  wire [63:0] cause; // @[CSR.scala 637:8]
  wire [7:0] cause_lsbs; // @[CSR.scala 639:25]
  wire  _T_1146; // @[CSR.scala 640:53]
  wire  causeIsDebugInt; // @[CSR.scala 640:39]
  wire  _T_1158; // @[CSR.scala 643:60]
  wire  causeIsDebugTrigger; // @[CSR.scala 641:44]
  wire  _T_1159; // @[CSR.scala 643:79]
  wire  _T_1152; // @[CSR.scala 642:42]
  reg  reg_dcsr_ebreakm; // @[CSR.scala 320:21]
  reg [31:0] _RAND_16;
  reg  reg_dcsr_ebreaks; // @[CSR.scala 320:21]
  reg [31:0] _RAND_17;
  reg  reg_dcsr_ebreaku; // @[CSR.scala 320:21]
  reg [31:0] _RAND_18;
  wire [3:0] _T_1155; // @[Cat.scala 29:58]
  wire [3:0] _T_1156; // @[CSR.scala 642:134]
  wire  causeIsDebugBreak; // @[CSR.scala 642:56]
  wire  _T_1160; // @[CSR.scala 643:102]
  reg  reg_debug; // @[CSR.scala 361:22]
  reg [31:0] _RAND_19;
  wire  trapToDebug; // @[CSR.scala 643:123]
  wire [1:0] _GEN_42; // @[CSR.scala 690:25]
  wire  _T_1163; // @[CSR.scala 645:59]
  reg [63:0] reg_mideleg; // @[CSR.scala 372:18]
  reg [63:0] _RAND_20;
  wire [63:0] read_mideleg; // @[CSR.scala 373:36]
  wire [63:0] _T_1166; // @[CSR.scala 645:102]
  reg [63:0] reg_medeleg; // @[CSR.scala 376:18]
  reg [63:0] _RAND_21;
  wire [63:0] read_medeleg; // @[CSR.scala 377:36]
  wire [63:0] _T_1168; // @[CSR.scala 645:128]
  wire  _T_1170; // @[CSR.scala 645:74]
  wire  delegate; // @[CSR.scala 645:68]
  wire [1:0] _GEN_50; // @[CSR.scala 697:27]
  wire [1:0] _GEN_61; // @[CSR.scala 689:24]
  wire [1:0] _GEN_79; // @[CSR.scala 688:20]
  wire [1:0] new_prv; // @[CSR.scala 738:19]
  wire  _T_1; // @[CSR.scala 1073:35]
  reg [2:0] reg_dcsr_cause; // @[CSR.scala 320:21]
  reg [31:0] _RAND_22;
  reg  reg_dcsr_step; // @[CSR.scala 320:21]
  reg [31:0] _RAND_23;
  reg [39:0] reg_dpc; // @[CSR.scala 362:20]
  reg [63:0] _RAND_24;
  reg [63:0] reg_dscratch; // @[CSR.scala 363:25]
  reg [63:0] _RAND_25;
  reg  reg_bp_0_control_dmode; // @[CSR.scala 367:19]
  reg [31:0] _RAND_26;
  reg  reg_bp_0_control_action; // @[CSR.scala 367:19]
  reg [31:0] _RAND_27;
  reg [1:0] reg_bp_0_control_tmatch; // @[CSR.scala 367:19]
  reg [31:0] _RAND_28;
  reg  reg_bp_0_control_m; // @[CSR.scala 367:19]
  reg [31:0] _RAND_29;
  reg  reg_bp_0_control_s; // @[CSR.scala 367:19]
  reg [31:0] _RAND_30;
  reg  reg_bp_0_control_u; // @[CSR.scala 367:19]
  reg [31:0] _RAND_31;
  reg  reg_bp_0_control_x; // @[CSR.scala 367:19]
  reg [31:0] _RAND_32;
  reg  reg_bp_0_control_w; // @[CSR.scala 367:19]
  reg [31:0] _RAND_33;
  reg  reg_bp_0_control_r; // @[CSR.scala 367:19]
  reg [31:0] _RAND_34;
  reg [38:0] reg_bp_0_address; // @[CSR.scala 367:19]
  reg [63:0] _RAND_35;
  reg  reg_pmp_0_cfg_l; // @[CSR.scala 368:20]
  reg [31:0] _RAND_36;
  reg [1:0] reg_pmp_0_cfg_a; // @[CSR.scala 368:20]
  reg [31:0] _RAND_37;
  reg  reg_pmp_0_cfg_x; // @[CSR.scala 368:20]
  reg [31:0] _RAND_38;
  reg  reg_pmp_0_cfg_w; // @[CSR.scala 368:20]
  reg [31:0] _RAND_39;
  reg  reg_pmp_0_cfg_r; // @[CSR.scala 368:20]
  reg [31:0] _RAND_40;
  reg [29:0] reg_pmp_0_addr; // @[CSR.scala 368:20]
  reg [31:0] _RAND_41;
  reg  reg_pmp_1_cfg_l; // @[CSR.scala 368:20]
  reg [31:0] _RAND_42;
  reg [1:0] reg_pmp_1_cfg_a; // @[CSR.scala 368:20]
  reg [31:0] _RAND_43;
  reg  reg_pmp_1_cfg_x; // @[CSR.scala 368:20]
  reg [31:0] _RAND_44;
  reg  reg_pmp_1_cfg_w; // @[CSR.scala 368:20]
  reg [31:0] _RAND_45;
  reg  reg_pmp_1_cfg_r; // @[CSR.scala 368:20]
  reg [31:0] _RAND_46;
  reg [29:0] reg_pmp_1_addr; // @[CSR.scala 368:20]
  reg [31:0] _RAND_47;
  reg  reg_pmp_2_cfg_l; // @[CSR.scala 368:20]
  reg [31:0] _RAND_48;
  reg [1:0] reg_pmp_2_cfg_a; // @[CSR.scala 368:20]
  reg [31:0] _RAND_49;
  reg  reg_pmp_2_cfg_x; // @[CSR.scala 368:20]
  reg [31:0] _RAND_50;
  reg  reg_pmp_2_cfg_w; // @[CSR.scala 368:20]
  reg [31:0] _RAND_51;
  reg  reg_pmp_2_cfg_r; // @[CSR.scala 368:20]
  reg [31:0] _RAND_52;
  reg [29:0] reg_pmp_2_addr; // @[CSR.scala 368:20]
  reg [31:0] _RAND_53;
  reg  reg_pmp_3_cfg_l; // @[CSR.scala 368:20]
  reg [31:0] _RAND_54;
  reg [1:0] reg_pmp_3_cfg_a; // @[CSR.scala 368:20]
  reg [31:0] _RAND_55;
  reg  reg_pmp_3_cfg_x; // @[CSR.scala 368:20]
  reg [31:0] _RAND_56;
  reg  reg_pmp_3_cfg_w; // @[CSR.scala 368:20]
  reg [31:0] _RAND_57;
  reg  reg_pmp_3_cfg_r; // @[CSR.scala 368:20]
  reg [31:0] _RAND_58;
  reg [29:0] reg_pmp_3_addr; // @[CSR.scala 368:20]
  reg [31:0] _RAND_59;
  reg  reg_pmp_4_cfg_l; // @[CSR.scala 368:20]
  reg [31:0] _RAND_60;
  reg [1:0] reg_pmp_4_cfg_a; // @[CSR.scala 368:20]
  reg [31:0] _RAND_61;
  reg  reg_pmp_4_cfg_x; // @[CSR.scala 368:20]
  reg [31:0] _RAND_62;
  reg  reg_pmp_4_cfg_w; // @[CSR.scala 368:20]
  reg [31:0] _RAND_63;
  reg  reg_pmp_4_cfg_r; // @[CSR.scala 368:20]
  reg [31:0] _RAND_64;
  reg [29:0] reg_pmp_4_addr; // @[CSR.scala 368:20]
  reg [31:0] _RAND_65;
  reg  reg_pmp_5_cfg_l; // @[CSR.scala 368:20]
  reg [31:0] _RAND_66;
  reg [1:0] reg_pmp_5_cfg_a; // @[CSR.scala 368:20]
  reg [31:0] _RAND_67;
  reg  reg_pmp_5_cfg_x; // @[CSR.scala 368:20]
  reg [31:0] _RAND_68;
  reg  reg_pmp_5_cfg_w; // @[CSR.scala 368:20]
  reg [31:0] _RAND_69;
  reg  reg_pmp_5_cfg_r; // @[CSR.scala 368:20]
  reg [31:0] _RAND_70;
  reg [29:0] reg_pmp_5_addr; // @[CSR.scala 368:20]
  reg [31:0] _RAND_71;
  reg  reg_pmp_6_cfg_l; // @[CSR.scala 368:20]
  reg [31:0] _RAND_72;
  reg [1:0] reg_pmp_6_cfg_a; // @[CSR.scala 368:20]
  reg [31:0] _RAND_73;
  reg  reg_pmp_6_cfg_x; // @[CSR.scala 368:20]
  reg [31:0] _RAND_74;
  reg  reg_pmp_6_cfg_w; // @[CSR.scala 368:20]
  reg [31:0] _RAND_75;
  reg  reg_pmp_6_cfg_r; // @[CSR.scala 368:20]
  reg [31:0] _RAND_76;
  reg [29:0] reg_pmp_6_addr; // @[CSR.scala 368:20]
  reg [31:0] _RAND_77;
  reg  reg_pmp_7_cfg_l; // @[CSR.scala 368:20]
  reg [31:0] _RAND_78;
  reg [1:0] reg_pmp_7_cfg_a; // @[CSR.scala 368:20]
  reg [31:0] _RAND_79;
  reg  reg_pmp_7_cfg_x; // @[CSR.scala 368:20]
  reg [31:0] _RAND_80;
  reg  reg_pmp_7_cfg_w; // @[CSR.scala 368:20]
  reg [31:0] _RAND_81;
  reg  reg_pmp_7_cfg_r; // @[CSR.scala 368:20]
  reg [31:0] _RAND_82;
  reg [29:0] reg_pmp_7_addr; // @[CSR.scala 368:20]
  reg [31:0] _RAND_83;
  reg [63:0] reg_mie; // @[CSR.scala 370:20]
  reg [63:0] _RAND_84;
  reg  reg_mip_seip; // @[CSR.scala 379:20]
  reg [31:0] _RAND_85;
  reg  reg_mip_stip; // @[CSR.scala 379:20]
  reg [31:0] _RAND_86;
  reg  reg_mip_ssip; // @[CSR.scala 379:20]
  reg [31:0] _RAND_87;
  reg [39:0] reg_mepc; // @[CSR.scala 380:21]
  reg [63:0] _RAND_88;
  reg [63:0] reg_mcause; // @[CSR.scala 381:27]
  reg [63:0] _RAND_89;
  reg [39:0] reg_mtval; // @[CSR.scala 382:22]
  reg [63:0] _RAND_90;
  reg [63:0] reg_mscratch; // @[CSR.scala 383:25]
  reg [63:0] _RAND_91;
  reg [31:0] reg_mtvec; // @[CSR.scala 386:27]
  reg [31:0] _RAND_92;
  reg [31:0] reg_mcounteren; // @[CSR.scala 392:18]
  reg [31:0] _RAND_93;
  wire [31:0] read_mcounteren; // @[CSR.scala 393:30]
  reg [31:0] reg_scounteren; // @[CSR.scala 396:18]
  reg [31:0] _RAND_94;
  wire [31:0] read_scounteren; // @[CSR.scala 397:36]
  reg [39:0] reg_sepc; // @[CSR.scala 400:21]
  reg [63:0] _RAND_95;
  reg [63:0] reg_scause; // @[CSR.scala 401:23]
  reg [63:0] _RAND_96;
  reg [39:0] reg_stval; // @[CSR.scala 402:22]
  reg [63:0] _RAND_97;
  reg [63:0] reg_sscratch; // @[CSR.scala 403:25]
  reg [63:0] _RAND_98;
  reg [38:0] reg_stvec; // @[CSR.scala 404:22]
  reg [63:0] _RAND_99;
  reg [3:0] reg_satp_mode; // @[CSR.scala 405:21]
  reg [31:0] _RAND_100;
  reg [43:0] reg_satp_ppn; // @[CSR.scala 405:21]
  reg [63:0] _RAND_101;
  reg  reg_wfi; // @[CSR.scala 406:50]
  reg [31:0] _RAND_102;
  reg [4:0] reg_fflags; // @[CSR.scala 408:23]
  reg [31:0] _RAND_103;
  reg [2:0] reg_frm; // @[CSR.scala 409:20]
  reg [31:0] _RAND_104;
  reg [5:0] _T_39; // @[Counters.scala 46:37]
  reg [31:0] _RAND_105;
  wire [5:0] _GEN_491; // @[Counters.scala 47:33]
  wire [6:0] _T_40; // @[Counters.scala 47:33]
  reg [57:0] _T_41; // @[Counters.scala 51:27]
  reg [63:0] _RAND_106;
  wire [57:0] _T_44; // @[Counters.scala 52:43]
  wire [63:0] _T_45; // @[Cat.scala 29:58]
  reg [5:0] _T_47; // @[Counters.scala 46:37]
  reg [31:0] _RAND_107;
  wire [5:0] _GEN_492; // @[Counters.scala 47:33]
  wire [6:0] _T_48; // @[Counters.scala 47:33]
  reg [57:0] _T_49; // @[Counters.scala 51:27]
  reg [63:0] _RAND_108;
  wire [57:0] _T_52; // @[Counters.scala 52:43]
  wire [63:0] _T_53; // @[Cat.scala 29:58]
  wire  mip_seip; // @[CSR.scala 427:57]
  wire [7:0] _T_61; // @[CSR.scala 429:22]
  wire [15:0] _T_69; // @[CSR.scala 429:22]
  wire [15:0] read_mip; // @[CSR.scala 429:29]
  wire [63:0] _GEN_493; // @[CSR.scala 432:56]
  wire [63:0] pending_interrupts; // @[CSR.scala 432:56]
  wire [14:0] d_interrupts; // @[CSR.scala 433:42]
  wire  _T_72; // @[CSR.scala 434:51]
  wire [63:0] _T_74; // @[CSR.scala 434:93]
  wire [63:0] m_interrupts; // @[CSR.scala 434:25]
  wire  _T_76; // @[CSR.scala 435:42]
  wire  _T_77; // @[CSR.scala 435:70]
  wire  _T_78; // @[CSR.scala 435:80]
  wire  _T_79; // @[CSR.scala 435:50]
  wire [63:0] _T_80; // @[CSR.scala 435:120]
  wire [63:0] s_interrupts; // @[CSR.scala 435:25]
  wire  _T_119; // @[CSR.scala 1063:90]
  wire  _T_120; // @[CSR.scala 1063:90]
  wire  _T_121; // @[CSR.scala 1063:90]
  wire  _T_122; // @[CSR.scala 1063:90]
  wire  _T_123; // @[CSR.scala 1063:90]
  wire  _T_124; // @[CSR.scala 1063:90]
  wire  _T_125; // @[CSR.scala 1063:90]
  wire  _T_126; // @[CSR.scala 1063:90]
  wire  _T_127; // @[CSR.scala 1063:90]
  wire  _T_128; // @[CSR.scala 1063:90]
  wire  _T_129; // @[CSR.scala 1063:90]
  wire  _T_130; // @[CSR.scala 1063:90]
  wire  _T_131; // @[CSR.scala 1063:90]
  wire  _T_132; // @[CSR.scala 1063:90]
  wire  _T_133; // @[CSR.scala 1063:90]
  wire  _T_134; // @[CSR.scala 1063:90]
  wire  _T_135; // @[CSR.scala 1063:90]
  wire  _T_136; // @[CSR.scala 1063:90]
  wire  _T_137; // @[CSR.scala 1063:90]
  wire  _T_138; // @[CSR.scala 1063:90]
  wire  _T_139; // @[CSR.scala 1063:90]
  wire  _T_140; // @[CSR.scala 1063:90]
  wire  _T_141; // @[CSR.scala 1063:90]
  wire  _T_142; // @[CSR.scala 1063:90]
  wire  _T_143; // @[CSR.scala 1063:90]
  wire  _T_144; // @[CSR.scala 1063:90]
  wire  _T_145; // @[CSR.scala 1063:90]
  wire  _T_146; // @[CSR.scala 1063:90]
  wire  _T_147; // @[CSR.scala 1063:90]
  wire  _T_148; // @[CSR.scala 1063:90]
  wire  _T_149; // @[CSR.scala 1063:90]
  wire  _T_150; // @[CSR.scala 1063:90]
  wire  _T_151; // @[CSR.scala 1063:90]
  wire  _T_152; // @[CSR.scala 1063:90]
  wire  _T_153; // @[CSR.scala 1063:90]
  wire  _T_154; // @[CSR.scala 1063:90]
  wire  anyInterrupt; // @[CSR.scala 1063:90]
  wire [2:0] _T_193; // @[Mux.scala 47:69]
  wire [3:0] _T_194; // @[Mux.scala 47:69]
  wire [3:0] _T_195; // @[Mux.scala 47:69]
  wire [3:0] _T_196; // @[Mux.scala 47:69]
  wire [3:0] _T_197; // @[Mux.scala 47:69]
  wire [3:0] _T_198; // @[Mux.scala 47:69]
  wire [3:0] _T_199; // @[Mux.scala 47:69]
  wire [3:0] _T_200; // @[Mux.scala 47:69]
  wire [3:0] _T_201; // @[Mux.scala 47:69]
  wire [3:0] _T_202; // @[Mux.scala 47:69]
  wire [3:0] _T_203; // @[Mux.scala 47:69]
  wire [3:0] _T_204; // @[Mux.scala 47:69]
  wire [3:0] _T_205; // @[Mux.scala 47:69]
  wire [3:0] _T_206; // @[Mux.scala 47:69]
  wire [3:0] _T_207; // @[Mux.scala 47:69]
  wire [3:0] _T_208; // @[Mux.scala 47:69]
  wire [3:0] _T_209; // @[Mux.scala 47:69]
  wire [3:0] _T_210; // @[Mux.scala 47:69]
  wire [3:0] _T_211; // @[Mux.scala 47:69]
  wire [3:0] _T_212; // @[Mux.scala 47:69]
  wire [3:0] _T_213; // @[Mux.scala 47:69]
  wire [3:0] _T_214; // @[Mux.scala 47:69]
  wire [3:0] _T_215; // @[Mux.scala 47:69]
  wire [3:0] _T_216; // @[Mux.scala 47:69]
  wire [3:0] _T_217; // @[Mux.scala 47:69]
  wire [3:0] _T_218; // @[Mux.scala 47:69]
  wire [3:0] _T_219; // @[Mux.scala 47:69]
  wire [3:0] _T_220; // @[Mux.scala 47:69]
  wire [3:0] _T_221; // @[Mux.scala 47:69]
  wire [3:0] _T_222; // @[Mux.scala 47:69]
  wire [3:0] _T_223; // @[Mux.scala 47:69]
  wire [3:0] _T_224; // @[Mux.scala 47:69]
  wire [3:0] _T_225; // @[Mux.scala 47:69]
  wire [3:0] _T_226; // @[Mux.scala 47:69]
  wire [3:0] _T_227; // @[Mux.scala 47:69]
  wire [3:0] _T_228; // @[Mux.scala 47:69]
  wire [3:0] whichInterrupt; // @[Mux.scala 47:69]
  wire [63:0] _GEN_494; // @[CSR.scala 438:43]
  wire  _T_231; // @[CSR.scala 439:33]
  wire  _T_232; // @[CSR.scala 439:51]
  wire  _T_233; // @[CSR.scala 439:88]
  wire [30:0] _T_238; // @[Cat.scala 29:58]
  wire [30:0] _T_241; // @[PMP.scala 60:23]
  wire [30:0] _T_243; // @[PMP.scala 60:14]
  wire [32:0] _T_244; // @[Cat.scala 29:58]
  wire [30:0] _T_247; // @[Cat.scala 29:58]
  wire [30:0] _T_250; // @[PMP.scala 60:23]
  wire [30:0] _T_252; // @[PMP.scala 60:14]
  wire [32:0] _T_253; // @[Cat.scala 29:58]
  wire [30:0] _T_256; // @[Cat.scala 29:58]
  wire [30:0] _T_259; // @[PMP.scala 60:23]
  wire [30:0] _T_261; // @[PMP.scala 60:14]
  wire [32:0] _T_262; // @[Cat.scala 29:58]
  wire [30:0] _T_265; // @[Cat.scala 29:58]
  wire [30:0] _T_268; // @[PMP.scala 60:23]
  wire [30:0] _T_270; // @[PMP.scala 60:14]
  wire [32:0] _T_271; // @[Cat.scala 29:58]
  wire [30:0] _T_274; // @[Cat.scala 29:58]
  wire [30:0] _T_277; // @[PMP.scala 60:23]
  wire [30:0] _T_279; // @[PMP.scala 60:14]
  wire [32:0] _T_280; // @[Cat.scala 29:58]
  wire [30:0] _T_283; // @[Cat.scala 29:58]
  wire [30:0] _T_286; // @[PMP.scala 60:23]
  wire [30:0] _T_288; // @[PMP.scala 60:14]
  wire [32:0] _T_289; // @[Cat.scala 29:58]
  wire [30:0] _T_292; // @[Cat.scala 29:58]
  wire [30:0] _T_295; // @[PMP.scala 60:23]
  wire [30:0] _T_297; // @[PMP.scala 60:14]
  wire [32:0] _T_298; // @[Cat.scala 29:58]
  wire [30:0] _T_301; // @[Cat.scala 29:58]
  wire [30:0] _T_304; // @[PMP.scala 60:23]
  wire [30:0] _T_306; // @[PMP.scala 60:14]
  wire [32:0] _T_307; // @[Cat.scala 29:58]
  reg [63:0] reg_misa; // @[CSR.scala 457:21]
  reg [63:0] _RAND_109;
  wire [6:0] _T_313; // @[CSR.scala 458:38]
  wire [18:0] _T_321; // @[CSR.scala 458:38]
  wire [16:0] _T_328; // @[CSR.scala 458:38]
  wire [102:0] _T_337; // @[CSR.scala 458:38]
  wire [63:0] read_mstatus; // @[CSR.scala 458:40]
  wire [7:0] _T_339; // @[CSR.scala 1092:39]
  wire [31:0] _T_341; // @[package.scala 154:41]
  wire [31:0] _T_343; // @[package.scala 154:35]
  wire [63:0] read_mtvec; // @[Cat.scala 29:58]
  wire [7:0] _T_345; // @[CSR.scala 1092:39]
  wire [38:0] _T_347; // @[package.scala 154:41]
  wire [38:0] _T_349; // @[package.scala 154:35]
  wire [24:0] _T_352; // @[Bitwise.scala 72:12]
  wire [63:0] read_stvec; // @[Cat.scala 29:58]
  wire [6:0] _T_358; // @[CSR.scala 464:48]
  wire [63:0] _T_366; // @[CSR.scala 464:48]
  wire [24:0] _T_369; // @[Bitwise.scala 72:12]
  wire [63:0] _T_370; // @[Cat.scala 29:58]
  wire [1:0] _T_373; // @[CSR.scala 1091:36]
  wire [39:0] _GEN_495; // @[CSR.scala 1091:31]
  wire [39:0] _T_374; // @[CSR.scala 1091:31]
  wire  _T_376; // @[package.scala 112:38]
  wire [23:0] _T_378; // @[Bitwise.scala 72:12]
  wire [63:0] _T_379; // @[Cat.scala 29:58]
  wire [23:0] _T_382; // @[Bitwise.scala 72:12]
  wire [63:0] _T_383; // @[Cat.scala 29:58]
  wire [11:0] _T_389; // @[CSR.scala 478:27]
  wire [31:0] _T_396; // @[CSR.scala 478:27]
  wire [39:0] _T_400; // @[CSR.scala 1091:31]
  wire  _T_402; // @[package.scala 112:38]
  wire [23:0] _T_404; // @[Bitwise.scala 72:12]
  wire [63:0] _T_405; // @[Cat.scala 29:58]
  wire [7:0] read_fcsr; // @[Cat.scala 29:58]
  wire [63:0] _T_406; // @[CSR.scala 534:28]
  wire [63:0] _T_407; // @[CSR.scala 535:29]
  wire [6:0] _T_415; // @[CSR.scala 549:57]
  wire [18:0] _T_423; // @[CSR.scala 549:57]
  wire [16:0] _T_430; // @[CSR.scala 549:57]
  wire [102:0] _T_439; // @[CSR.scala 549:57]
  wire [23:0] _T_443; // @[Bitwise.scala 72:12]
  wire [63:0] _T_444; // @[Cat.scala 29:58]
  wire [63:0] _T_446; // @[CSR.scala 555:43]
  wire [39:0] _T_450; // @[CSR.scala 1091:31]
  wire  _T_452; // @[package.scala 112:38]
  wire [23:0] _T_454; // @[Bitwise.scala 72:12]
  wire [63:0] _T_455; // @[Cat.scala 29:58]
  wire [7:0] _T_461; // @[package.scala 36:38]
  wire [7:0] _T_471; // @[package.scala 36:38]
  wire [7:0] _T_481; // @[package.scala 36:38]
  wire [7:0] _T_491; // @[package.scala 36:38]
  wire [15:0] _T_497; // @[Cat.scala 29:58]
  wire [31:0] _T_499; // @[Cat.scala 29:58]
  wire [15:0] _T_500; // @[Cat.scala 29:58]
  wire [63:0] _T_503; // @[Cat.scala 29:58]
  reg [63:0] reg_custom_0; // @[CSR.scala 578:43]
  reg [63:0] _RAND_110;
  wire  _T_552; // @[CSR.scala 586:73]
  wire  _T_553; // @[CSR.scala 586:73]
  wire  _T_554; // @[CSR.scala 586:73]
  wire  _T_555; // @[CSR.scala 586:73]
  wire  _T_556; // @[CSR.scala 586:73]
  wire  _T_557; // @[CSR.scala 586:73]
  wire  _T_558; // @[CSR.scala 586:73]
  wire  _T_559; // @[CSR.scala 586:73]
  wire  _T_560; // @[CSR.scala 586:73]
  wire  _T_561; // @[CSR.scala 586:73]
  wire  _T_562; // @[CSR.scala 586:73]
  wire  _T_563; // @[CSR.scala 586:73]
  wire  _T_564; // @[CSR.scala 586:73]
  wire  _T_565; // @[CSR.scala 586:73]
  wire  _T_566; // @[CSR.scala 586:73]
  wire  _T_567; // @[CSR.scala 586:73]
  wire  _T_568; // @[CSR.scala 586:73]
  wire  _T_569; // @[CSR.scala 586:73]
  wire  _T_570; // @[CSR.scala 586:73]
  wire  _T_571; // @[CSR.scala 586:73]
  wire  _T_659; // @[CSR.scala 586:73]
  wire  _T_660; // @[CSR.scala 586:73]
  wire  _T_661; // @[CSR.scala 586:73]
  wire  _T_662; // @[CSR.scala 586:73]
  wire  _T_663; // @[CSR.scala 586:73]
  wire  _T_664; // @[CSR.scala 586:73]
  wire  _T_665; // @[CSR.scala 586:73]
  wire  _T_666; // @[CSR.scala 586:73]
  wire  _T_667; // @[CSR.scala 586:73]
  wire  _T_668; // @[CSR.scala 586:73]
  wire  _T_669; // @[CSR.scala 586:73]
  wire  _T_670; // @[CSR.scala 586:73]
  wire  _T_671; // @[CSR.scala 586:73]
  wire  _T_672; // @[CSR.scala 586:73]
  wire  _T_673; // @[CSR.scala 586:73]
  wire  _T_674; // @[CSR.scala 586:73]
  wire  _T_676; // @[CSR.scala 586:73]
  wire  _T_677; // @[CSR.scala 586:73]
  wire  _T_678; // @[CSR.scala 586:73]
  wire  _T_679; // @[CSR.scala 586:73]
  wire  _T_680; // @[CSR.scala 586:73]
  wire  _T_681; // @[CSR.scala 586:73]
  wire  _T_682; // @[CSR.scala 586:73]
  wire  _T_683; // @[CSR.scala 586:73]
  wire  _T_692; // @[CSR.scala 586:73]
  wire  _T_693; // @[CSR.scala 586:73]
  wire  _T_695; // @[CSR.scala 586:73]
  wire [63:0] _T_697; // @[CSR.scala 1069:9]
  wire [63:0] _T_698; // @[CSR.scala 1069:34]
  wire  _T_700; // @[CSR.scala 1069:59]
  wire [63:0] _T_701; // @[CSR.scala 1069:49]
  wire [63:0] wdata; // @[CSR.scala 1069:43]
  wire [31:0] _T_716; // @[Decode.scala 14:65]
  wire  _T_717; // @[Decode.scala 14:121]
  wire [31:0] _T_719; // @[Decode.scala 14:65]
  wire  _T_720; // @[Decode.scala 14:121]
  wire  insn_cease; // @[CSR.scala 601:95]
  wire  insn_wfi; // @[CSR.scala 601:95]
  wire [31:0] _T_731; // @[CSR.scala 608:30]
  wire [31:0] _T_738; // @[Decode.scala 14:65]
  wire  _T_739; // @[Decode.scala 14:121]
  wire [31:0] _T_740; // @[Decode.scala 14:65]
  wire  _T_741; // @[Decode.scala 14:121]
  wire  _T_743; // @[Decode.scala 15:30]
  wire [31:0] _T_747; // @[Decode.scala 14:65]
  wire  _T_748; // @[Decode.scala 14:121]
  wire [31:0] _T_750; // @[Decode.scala 14:65]
  wire  _T_751; // @[Decode.scala 14:121]
  wire  _T_759; // @[CSR.scala 610:63]
  wire  _T_762; // @[CSR.scala 610:71]
  wire  _T_766; // @[CSR.scala 611:70]
  wire  _T_770; // @[CSR.scala 612:72]
  wire [31:0] _T_773; // @[CSR.scala 614:68]
  wire  _T_775; // @[CSR.scala 614:50]
  wire  _T_776; // @[CSR.scala 615:44]
  wire [31:0] _T_778; // @[CSR.scala 615:71]
  wire  _T_780; // @[CSR.scala 615:53]
  wire  _T_781; // @[CSR.scala 614:84]
  wire  _T_782; // @[CSR.scala 616:39]
  wire [11:0] _T_790; // @[Decode.scala 14:65]
  wire  _T_799; // @[CSR.scala 620:44]
  wire  _T_800; // @[CSR.scala 604:99]
  wire  _T_801; // @[CSR.scala 604:99]
  wire  _T_802; // @[CSR.scala 604:99]
  wire  _T_803; // @[CSR.scala 604:99]
  wire  _T_804; // @[CSR.scala 604:99]
  wire  _T_805; // @[CSR.scala 604:99]
  wire  _T_806; // @[CSR.scala 604:99]
  wire  _T_807; // @[CSR.scala 604:99]
  wire  _T_808; // @[CSR.scala 604:99]
  wire  _T_809; // @[CSR.scala 604:99]
  wire  _T_810; // @[CSR.scala 604:99]
  wire  _T_811; // @[CSR.scala 604:99]
  wire  _T_812; // @[CSR.scala 604:99]
  wire  _T_813; // @[CSR.scala 604:99]
  wire  _T_814; // @[CSR.scala 604:99]
  wire  _T_815; // @[CSR.scala 604:99]
  wire  _T_816; // @[CSR.scala 604:99]
  wire  _T_817; // @[CSR.scala 604:99]
  wire  _T_818; // @[CSR.scala 604:99]
  wire  _T_819; // @[CSR.scala 604:99]
  wire  _T_820; // @[CSR.scala 604:99]
  wire  _T_821; // @[CSR.scala 604:99]
  wire  _T_822; // @[CSR.scala 604:99]
  wire  _T_823; // @[CSR.scala 604:99]
  wire  _T_824; // @[CSR.scala 604:99]
  wire  _T_825; // @[CSR.scala 604:99]
  wire  _T_826; // @[CSR.scala 604:99]
  wire  _T_827; // @[CSR.scala 604:99]
  wire  _T_828; // @[CSR.scala 604:99]
  wire  _T_829; // @[CSR.scala 604:99]
  wire  _T_830; // @[CSR.scala 604:99]
  wire  _T_831; // @[CSR.scala 604:99]
  wire  _T_832; // @[CSR.scala 604:99]
  wire  _T_833; // @[CSR.scala 604:99]
  wire  _T_834; // @[CSR.scala 604:99]
  wire  _T_835; // @[CSR.scala 604:99]
  wire  _T_836; // @[CSR.scala 604:99]
  wire  _T_837; // @[CSR.scala 604:99]
  wire  _T_838; // @[CSR.scala 604:99]
  wire  _T_839; // @[CSR.scala 604:99]
  wire  _T_840; // @[CSR.scala 604:99]
  wire  _T_841; // @[CSR.scala 604:99]
  wire  _T_842; // @[CSR.scala 604:99]
  wire  _T_843; // @[CSR.scala 604:99]
  wire  _T_844; // @[CSR.scala 604:99]
  wire  _T_845; // @[CSR.scala 604:99]
  wire  _T_846; // @[CSR.scala 604:99]
  wire  _T_847; // @[CSR.scala 604:99]
  wire  _T_848; // @[CSR.scala 604:99]
  wire  _T_849; // @[CSR.scala 604:99]
  wire  _T_850; // @[CSR.scala 604:99]
  wire  _T_851; // @[CSR.scala 604:99]
  wire  _T_852; // @[CSR.scala 604:99]
  wire  _T_853; // @[CSR.scala 604:99]
  wire  _T_854; // @[CSR.scala 604:99]
  wire  _T_855; // @[CSR.scala 604:99]
  wire  _T_856; // @[CSR.scala 604:99]
  wire  _T_857; // @[CSR.scala 604:99]
  wire  _T_858; // @[CSR.scala 604:99]
  wire  _T_859; // @[CSR.scala 604:99]
  wire  _T_860; // @[CSR.scala 604:99]
  wire  _T_861; // @[CSR.scala 604:99]
  wire  _T_862; // @[CSR.scala 604:99]
  wire  _T_863; // @[CSR.scala 604:99]
  wire  _T_864; // @[CSR.scala 604:99]
  wire  _T_865; // @[CSR.scala 604:99]
  wire  _T_866; // @[CSR.scala 604:99]
  wire  _T_867; // @[CSR.scala 604:99]
  wire  _T_868; // @[CSR.scala 604:99]
  wire  _T_869; // @[CSR.scala 604:99]
  wire  _T_870; // @[CSR.scala 604:99]
  wire  _T_871; // @[CSR.scala 604:99]
  wire  _T_872; // @[CSR.scala 604:99]
  wire  _T_873; // @[CSR.scala 604:99]
  wire  _T_874; // @[CSR.scala 604:99]
  wire  _T_875; // @[CSR.scala 604:99]
  wire  _T_876; // @[CSR.scala 604:99]
  wire  _T_877; // @[CSR.scala 604:99]
  wire  _T_878; // @[CSR.scala 604:99]
  wire  _T_879; // @[CSR.scala 604:99]
  wire  _T_880; // @[CSR.scala 604:99]
  wire  _T_881; // @[CSR.scala 604:99]
  wire  _T_882; // @[CSR.scala 604:99]
  wire  _T_883; // @[CSR.scala 604:99]
  wire  _T_884; // @[CSR.scala 604:99]
  wire  _T_885; // @[CSR.scala 604:99]
  wire  _T_886; // @[CSR.scala 604:99]
  wire  _T_887; // @[CSR.scala 604:99]
  wire  _T_888; // @[CSR.scala 604:99]
  wire  _T_889; // @[CSR.scala 604:99]
  wire  _T_890; // @[CSR.scala 604:99]
  wire  _T_891; // @[CSR.scala 604:99]
  wire  _T_892; // @[CSR.scala 604:99]
  wire  _T_893; // @[CSR.scala 604:99]
  wire  _T_894; // @[CSR.scala 604:99]
  wire  _T_895; // @[CSR.scala 604:99]
  wire  _T_896; // @[CSR.scala 604:99]
  wire  _T_897; // @[CSR.scala 604:99]
  wire  _T_898; // @[CSR.scala 604:99]
  wire  _T_899; // @[CSR.scala 604:99]
  wire  _T_900; // @[CSR.scala 604:99]
  wire  _T_901; // @[CSR.scala 604:99]
  wire  _T_902; // @[CSR.scala 604:99]
  wire  _T_903; // @[CSR.scala 604:99]
  wire  _T_904; // @[CSR.scala 604:99]
  wire  _T_905; // @[CSR.scala 604:99]
  wire  _T_906; // @[CSR.scala 604:99]
  wire  _T_907; // @[CSR.scala 604:99]
  wire  _T_908; // @[CSR.scala 604:99]
  wire  _T_909; // @[CSR.scala 604:99]
  wire  _T_910; // @[CSR.scala 604:99]
  wire  _T_911; // @[CSR.scala 604:99]
  wire  _T_912; // @[CSR.scala 604:99]
  wire  _T_913; // @[CSR.scala 604:99]
  wire  _T_914; // @[CSR.scala 604:99]
  wire  _T_915; // @[CSR.scala 604:99]
  wire  _T_916; // @[CSR.scala 604:99]
  wire  _T_917; // @[CSR.scala 604:99]
  wire  _T_918; // @[CSR.scala 604:99]
  wire  _T_919; // @[CSR.scala 604:99]
  wire  _T_920; // @[CSR.scala 604:99]
  wire  _T_921; // @[CSR.scala 604:99]
  wire  _T_922; // @[CSR.scala 604:99]
  wire  _T_923; // @[CSR.scala 604:99]
  wire  _T_924; // @[CSR.scala 604:99]
  wire  _T_925; // @[CSR.scala 604:99]
  wire  _T_926; // @[CSR.scala 604:99]
  wire  _T_927; // @[CSR.scala 604:99]
  wire  _T_928; // @[CSR.scala 604:99]
  wire  _T_929; // @[CSR.scala 604:99]
  wire  _T_930; // @[CSR.scala 604:99]
  wire  _T_931; // @[CSR.scala 604:99]
  wire  _T_932; // @[CSR.scala 604:99]
  wire  _T_933; // @[CSR.scala 604:99]
  wire  _T_934; // @[CSR.scala 604:99]
  wire  _T_935; // @[CSR.scala 604:99]
  wire  _T_936; // @[CSR.scala 604:99]
  wire  _T_937; // @[CSR.scala 604:99]
  wire  _T_938; // @[CSR.scala 604:99]
  wire  _T_939; // @[CSR.scala 604:99]
  wire  _T_940; // @[CSR.scala 604:99]
  wire  _T_941; // @[CSR.scala 604:99]
  wire  _T_942; // @[CSR.scala 604:99]
  wire  _T_943; // @[CSR.scala 604:99]
  wire  _T_944; // @[CSR.scala 604:99]
  wire  _T_945; // @[CSR.scala 604:115]
  wire  _T_946; // @[CSR.scala 604:115]
  wire  _T_947; // @[CSR.scala 604:115]
  wire  _T_948; // @[CSR.scala 604:115]
  wire  _T_949; // @[CSR.scala 604:115]
  wire  _T_950; // @[CSR.scala 604:115]
  wire  _T_951; // @[CSR.scala 604:115]
  wire  _T_952; // @[CSR.scala 604:115]
  wire  _T_953; // @[CSR.scala 604:115]
  wire  _T_954; // @[CSR.scala 604:115]
  wire  _T_955; // @[CSR.scala 604:115]
  wire  _T_956; // @[CSR.scala 604:115]
  wire  _T_957; // @[CSR.scala 604:115]
  wire  _T_958; // @[CSR.scala 604:115]
  wire  _T_959; // @[CSR.scala 604:115]
  wire  _T_960; // @[CSR.scala 604:115]
  wire  _T_961; // @[CSR.scala 604:115]
  wire  _T_962; // @[CSR.scala 604:115]
  wire  _T_963; // @[CSR.scala 604:115]
  wire  _T_964; // @[CSR.scala 604:115]
  wire  _T_965; // @[CSR.scala 604:115]
  wire  _T_966; // @[CSR.scala 604:115]
  wire  _T_967; // @[CSR.scala 604:115]
  wire  _T_968; // @[CSR.scala 604:115]
  wire  _T_969; // @[CSR.scala 604:115]
  wire  _T_970; // @[CSR.scala 604:115]
  wire  _T_971; // @[CSR.scala 604:115]
  wire  _T_972; // @[CSR.scala 604:115]
  wire  _T_973; // @[CSR.scala 604:115]
  wire  _T_974; // @[CSR.scala 604:115]
  wire  _T_975; // @[CSR.scala 604:115]
  wire  _T_976; // @[CSR.scala 604:115]
  wire  _T_977; // @[CSR.scala 604:115]
  wire  _T_978; // @[CSR.scala 604:115]
  wire  _T_979; // @[CSR.scala 604:115]
  wire  _T_980; // @[CSR.scala 604:115]
  wire  _T_981; // @[CSR.scala 604:115]
  wire  _T_982; // @[CSR.scala 604:115]
  wire  _T_983; // @[CSR.scala 604:115]
  wire  _T_984; // @[CSR.scala 604:115]
  wire  _T_985; // @[CSR.scala 604:115]
  wire  _T_986; // @[CSR.scala 604:115]
  wire  _T_987; // @[CSR.scala 604:115]
  wire  _T_988; // @[CSR.scala 604:115]
  wire  _T_989; // @[CSR.scala 604:115]
  wire  _T_990; // @[CSR.scala 604:115]
  wire  _T_991; // @[CSR.scala 604:115]
  wire  _T_992; // @[CSR.scala 604:115]
  wire  _T_993; // @[CSR.scala 604:115]
  wire  _T_994; // @[CSR.scala 604:115]
  wire  _T_995; // @[CSR.scala 604:115]
  wire  _T_996; // @[CSR.scala 604:115]
  wire  _T_997; // @[CSR.scala 604:115]
  wire  _T_998; // @[CSR.scala 604:115]
  wire  _T_999; // @[CSR.scala 604:115]
  wire  _T_1000; // @[CSR.scala 604:115]
  wire  _T_1001; // @[CSR.scala 604:115]
  wire  _T_1002; // @[CSR.scala 604:115]
  wire  _T_1003; // @[CSR.scala 604:115]
  wire  _T_1004; // @[CSR.scala 604:115]
  wire  _T_1005; // @[CSR.scala 604:115]
  wire  _T_1006; // @[CSR.scala 604:115]
  wire  _T_1007; // @[CSR.scala 604:115]
  wire  _T_1008; // @[CSR.scala 604:115]
  wire  _T_1009; // @[CSR.scala 604:115]
  wire  _T_1010; // @[CSR.scala 604:115]
  wire  _T_1011; // @[CSR.scala 604:115]
  wire  _T_1012; // @[CSR.scala 604:115]
  wire  _T_1013; // @[CSR.scala 604:115]
  wire  _T_1014; // @[CSR.scala 604:115]
  wire  _T_1015; // @[CSR.scala 604:115]
  wire  _T_1016; // @[CSR.scala 604:115]
  wire  _T_1017; // @[CSR.scala 604:115]
  wire  _T_1018; // @[CSR.scala 604:115]
  wire  _T_1019; // @[CSR.scala 604:115]
  wire  _T_1020; // @[CSR.scala 604:115]
  wire  _T_1021; // @[CSR.scala 604:115]
  wire  _T_1022; // @[CSR.scala 604:115]
  wire  _T_1023; // @[CSR.scala 604:115]
  wire  _T_1024; // @[CSR.scala 604:115]
  wire  _T_1025; // @[CSR.scala 604:115]
  wire  _T_1026; // @[CSR.scala 604:115]
  wire  _T_1027; // @[CSR.scala 604:115]
  wire  _T_1028; // @[CSR.scala 604:115]
  wire  _T_1029; // @[CSR.scala 604:115]
  wire  _T_1030; // @[CSR.scala 604:115]
  wire  _T_1031; // @[CSR.scala 604:115]
  wire  _T_1032; // @[CSR.scala 604:115]
  wire  _T_1033; // @[CSR.scala 604:115]
  wire  _T_1034; // @[CSR.scala 604:115]
  wire  _T_1035; // @[CSR.scala 604:115]
  wire  _T_1036; // @[CSR.scala 604:115]
  wire  _T_1037; // @[CSR.scala 604:115]
  wire  _T_1038; // @[CSR.scala 604:115]
  wire  _T_1039; // @[CSR.scala 604:115]
  wire  _T_1040; // @[CSR.scala 604:115]
  wire  _T_1041; // @[CSR.scala 604:115]
  wire  _T_1042; // @[CSR.scala 604:115]
  wire  _T_1043; // @[CSR.scala 604:115]
  wire  _T_1044; // @[CSR.scala 604:115]
  wire  _T_1045; // @[CSR.scala 604:115]
  wire  _T_1046; // @[CSR.scala 604:115]
  wire  _T_1047; // @[CSR.scala 604:115]
  wire  _T_1048; // @[CSR.scala 604:115]
  wire  _T_1049; // @[CSR.scala 604:115]
  wire  _T_1050; // @[CSR.scala 604:115]
  wire  _T_1051; // @[CSR.scala 604:115]
  wire  _T_1052; // @[CSR.scala 604:115]
  wire  _T_1053; // @[CSR.scala 604:115]
  wire  _T_1054; // @[CSR.scala 604:115]
  wire  _T_1055; // @[CSR.scala 604:115]
  wire  _T_1056; // @[CSR.scala 604:115]
  wire  _T_1057; // @[CSR.scala 604:115]
  wire  _T_1058; // @[CSR.scala 604:115]
  wire  _T_1059; // @[CSR.scala 604:115]
  wire  _T_1060; // @[CSR.scala 604:115]
  wire  _T_1061; // @[CSR.scala 604:115]
  wire  _T_1062; // @[CSR.scala 604:115]
  wire  _T_1063; // @[CSR.scala 604:115]
  wire  _T_1064; // @[CSR.scala 604:115]
  wire  _T_1065; // @[CSR.scala 604:115]
  wire  _T_1066; // @[CSR.scala 604:115]
  wire  _T_1067; // @[CSR.scala 604:115]
  wire  _T_1068; // @[CSR.scala 604:115]
  wire  _T_1069; // @[CSR.scala 604:115]
  wire  _T_1070; // @[CSR.scala 604:115]
  wire  _T_1071; // @[CSR.scala 604:115]
  wire  _T_1072; // @[CSR.scala 604:115]
  wire  _T_1073; // @[CSR.scala 604:115]
  wire  _T_1074; // @[CSR.scala 604:115]
  wire  _T_1075; // @[CSR.scala 604:115]
  wire  _T_1076; // @[CSR.scala 604:115]
  wire  _T_1077; // @[CSR.scala 604:115]
  wire  _T_1078; // @[CSR.scala 604:115]
  wire  _T_1079; // @[CSR.scala 604:115]
  wire  _T_1080; // @[CSR.scala 604:115]
  wire  _T_1081; // @[CSR.scala 604:115]
  wire  _T_1082; // @[CSR.scala 604:115]
  wire  _T_1083; // @[CSR.scala 604:115]
  wire  _T_1084; // @[CSR.scala 604:115]
  wire  _T_1085; // @[CSR.scala 604:115]
  wire  _T_1086; // @[CSR.scala 604:115]
  wire  _T_1087; // @[CSR.scala 604:115]
  wire  _T_1088; // @[CSR.scala 604:115]
  wire  _T_1090; // @[CSR.scala 620:62]
  wire  _T_1093; // @[CSR.scala 622:32]
  wire  _T_1094; // @[CSR.scala 621:32]
  wire  _T_1095; // @[package.scala 185:47]
  wire  _T_1096; // @[package.scala 185:60]
  wire  _T_1097; // @[package.scala 185:55]
  wire  _T_1098; // @[package.scala 185:47]
  wire  _T_1099; // @[package.scala 185:60]
  wire  _T_1100; // @[package.scala 185:55]
  wire  _T_1101; // @[CSR.scala 623:66]
  wire  _T_1103; // @[CSR.scala 623:130]
  wire  _T_1104; // @[CSR.scala 622:53]
  wire [11:0] _T_1105; // @[Decode.scala 14:65]
  wire  _T_1106; // @[Decode.scala 14:121]
  wire  _T_1110; // @[CSR.scala 624:42]
  wire  _T_1111; // @[CSR.scala 623:148]
  wire  _T_1114; // @[CSR.scala 626:21]
  wire  _T_1118; // @[CSR.scala 628:40]
  wire  _T_1119; // @[CSR.scala 628:71]
  wire  _T_1120; // @[CSR.scala 628:57]
  wire  _T_1121; // @[CSR.scala 628:99]
  wire  _T_1122; // @[CSR.scala 628:130]
  wire  _T_1123; // @[CSR.scala 628:116]
  wire  _T_1124; // @[CSR.scala 628:85]
  wire  _T_1129; // @[CSR.scala 630:14]
  wire  _T_1130; // @[CSR.scala 629:64]
  wire  _T_1132; // @[CSR.scala 631:14]
  wire  _T_1133; // @[CSR.scala 630:28]
  wire  _T_1135; // @[CSR.scala 632:14]
  wire  _T_1137; // @[CSR.scala 632:32]
  wire  _T_1138; // @[CSR.scala 631:29]
  wire  _T_1140; // @[CSR.scala 633:17]
  wire [11:0] _T_1162; // @[CSR.scala 644:37]
  wire [11:0] debugTVec; // @[CSR.scala 644:22]
  wire [63:0] _T_1171; // @[CSR.scala 652:19]
  wire [7:0] _T_1173; // @[CSR.scala 653:59]
  wire [63:0] _T_1175; // @[Cat.scala 29:58]
  wire  _T_1178; // @[CSR.scala 655:28]
  wire  _T_1180; // @[CSR.scala 655:94]
  wire  _T_1181; // @[CSR.scala 655:55]
  wire [63:0] _T_1183; // @[CSR.scala 656:56]
  wire [63:0] notDebugTVec; // @[CSR.scala 656:8]
  wire [63:0] tvec; // @[CSR.scala 658:17]
  wire  _T_1188; // @[CSR.scala 664:32]
  wire  _T_1189; // @[CSR.scala 664:53]
  wire  _T_1190; // @[CSR.scala 664:37]
  wire  _T_1191; // @[CSR.scala 664:74]
  wire  _T_1194; // @[CSR.scala 669:53]
  reg [1:0] _T_1196; // @[CSR.scala 669:24]
  reg [31:0] _RAND_111;
  wire [1:0] _T_1198; // @[Bitwise.scala 47:55]
  wire [1:0] _T_1200; // @[Bitwise.scala 47:55]
  wire [2:0] _T_1202; // @[Bitwise.scala 47:55]
  wire  _T_1204; // @[CSR.scala 674:79]
  wire  _T_1206; // @[CSR.scala 674:9]
  wire  _T_1209; // @[CSR.scala 676:18]
  wire  _T_1211; // @[CSR.scala 676:36]
  wire  _GEN_34; // @[CSR.scala 676:51]
  wire  _T_1212; // @[CSR.scala 677:28]
  wire  _T_1213; // @[CSR.scala 677:32]
  wire  _T_1214; // @[CSR.scala 677:55]
  wire  _T_1216; // @[CSR.scala 679:22]
  wire  _GEN_36; // @[CSR.scala 679:36]
  wire  _T_1226; // @[CSR.scala 682:29]
  wire  _T_1228; // @[CSR.scala 682:9]
  wire [39:0] _T_1231; // @[CSR.scala 1090:31]
  wire [39:0] epc; // @[CSR.scala 1090:26]
  wire [1:0] _T_1233; // @[CSR.scala 693:86]
  wire [1:0] _T_1234; // @[CSR.scala 693:56]
  wire  _GEN_38; // @[CSR.scala 690:25]
  wire [39:0] _GEN_39; // @[CSR.scala 690:25]
  wire [39:0] _GEN_43; // @[CSR.scala 697:27]
  wire  _GEN_47; // @[CSR.scala 697:27]
  wire [1:0] _GEN_48; // @[CSR.scala 697:27]
  wire [39:0] _GEN_51; // @[CSR.scala 697:27]
  wire  _GEN_54; // @[CSR.scala 697:27]
  wire [1:0] _GEN_55; // @[CSR.scala 697:27]
  wire  _GEN_56; // @[CSR.scala 697:27]
  wire [39:0] _GEN_58; // @[CSR.scala 689:24]
  wire [39:0] _GEN_62; // @[CSR.scala 689:24]
  wire  _GEN_66; // @[CSR.scala 689:24]
  wire [1:0] _GEN_67; // @[CSR.scala 689:24]
  wire [39:0] _GEN_69; // @[CSR.scala 689:24]
  wire  _GEN_72; // @[CSR.scala 689:24]
  wire [1:0] _GEN_73; // @[CSR.scala 689:24]
  wire  _GEN_74; // @[CSR.scala 689:24]
  wire [39:0] _GEN_76; // @[CSR.scala 688:20]
  wire [39:0] _GEN_80; // @[CSR.scala 688:20]
  wire  _GEN_84; // @[CSR.scala 688:20]
  wire [1:0] _GEN_85; // @[CSR.scala 688:20]
  wire [39:0] _GEN_87; // @[CSR.scala 688:20]
  wire  _GEN_90; // @[CSR.scala 688:20]
  wire [1:0] _GEN_91; // @[CSR.scala 688:20]
  wire  _GEN_92; // @[CSR.scala 688:20]
  wire [39:0] _GEN_95; // @[CSR.scala 745:53]
  wire  _GEN_100; // @[CSR.scala 739:52]
  wire [1:0] _GEN_101; // @[CSR.scala 739:52]
  wire [39:0] _GEN_103; // @[CSR.scala 739:52]
  wire [1:0] _GEN_110; // @[CSR.scala 738:19]
  wire [63:0] _GEN_112; // @[CSR.scala 738:19]
  reg  _T_1579; // @[Reg.scala 27:20]
  reg [31:0] _RAND_112;
  wire  _GEN_117; // @[Reg.scala 28:19]
  wire [63:0] _T_1581; // @[Mux.scala 27:72]
  wire [63:0] _T_1582; // @[Mux.scala 27:72]
  wire [63:0] _T_1583; // @[Mux.scala 27:72]
  wire [63:0] _T_1584; // @[Mux.scala 27:72]
  wire [63:0] _T_1585; // @[Mux.scala 27:72]
  wire [15:0] _T_1586; // @[Mux.scala 27:72]
  wire [63:0] _T_1587; // @[Mux.scala 27:72]
  wire [63:0] _T_1588; // @[Mux.scala 27:72]
  wire [63:0] _T_1589; // @[Mux.scala 27:72]
  wire [63:0] _T_1590; // @[Mux.scala 27:72]
  wire [63:0] _T_1591; // @[Mux.scala 27:72]
  wire  _T_1592; // @[Mux.scala 27:72]
  wire [31:0] _T_1593; // @[Mux.scala 27:72]
  wire [63:0] _T_1594; // @[Mux.scala 27:72]
  wire [63:0] _T_1595; // @[Mux.scala 27:72]
  wire [4:0] _T_1596; // @[Mux.scala 27:72]
  wire [2:0] _T_1597; // @[Mux.scala 27:72]
  wire [7:0] _T_1598; // @[Mux.scala 27:72]
  wire [63:0] _T_1599; // @[Mux.scala 27:72]
  wire [63:0] _T_1600; // @[Mux.scala 27:72]
  wire [31:0] _T_1688; // @[Mux.scala 27:72]
  wire [63:0] _T_1689; // @[Mux.scala 27:72]
  wire [63:0] _T_1690; // @[Mux.scala 27:72]
  wire [63:0] _T_1691; // @[Mux.scala 27:72]
  wire [63:0] _T_1692; // @[Mux.scala 27:72]
  wire [63:0] _T_1693; // @[Mux.scala 27:72]
  wire [63:0] _T_1694; // @[Mux.scala 27:72]
  wire [63:0] _T_1695; // @[Mux.scala 27:72]
  wire [63:0] _T_1696; // @[Mux.scala 27:72]
  wire [63:0] _T_1697; // @[Mux.scala 27:72]
  wire [63:0] _T_1698; // @[Mux.scala 27:72]
  wire [63:0] _T_1699; // @[Mux.scala 27:72]
  wire [31:0] _T_1700; // @[Mux.scala 27:72]
  wire [63:0] _T_1701; // @[Mux.scala 27:72]
  wire [63:0] _T_1702; // @[Mux.scala 27:72]
  wire [63:0] _T_1703; // @[Mux.scala 27:72]
  wire [29:0] _T_1705; // @[Mux.scala 27:72]
  wire [29:0] _T_1706; // @[Mux.scala 27:72]
  wire [29:0] _T_1707; // @[Mux.scala 27:72]
  wire [29:0] _T_1708; // @[Mux.scala 27:72]
  wire [29:0] _T_1709; // @[Mux.scala 27:72]
  wire [29:0] _T_1710; // @[Mux.scala 27:72]
  wire [29:0] _T_1711; // @[Mux.scala 27:72]
  wire [29:0] _T_1712; // @[Mux.scala 27:72]
  wire [63:0] _T_1721; // @[Mux.scala 27:72]
  wire [63:0] _T_1722; // @[Mux.scala 27:72]
  wire [63:0] _T_1724; // @[Mux.scala 27:72]
  wire [63:0] _T_1726; // @[Mux.scala 27:72]
  wire [63:0] _T_1727; // @[Mux.scala 27:72]
  wire [63:0] _T_1728; // @[Mux.scala 27:72]
  wire [63:0] _T_1729; // @[Mux.scala 27:72]
  wire [63:0] _GEN_502; // @[Mux.scala 27:72]
  wire [63:0] _T_1730; // @[Mux.scala 27:72]
  wire [63:0] _T_1731; // @[Mux.scala 27:72]
  wire [63:0] _T_1732; // @[Mux.scala 27:72]
  wire [63:0] _T_1733; // @[Mux.scala 27:72]
  wire [63:0] _T_1734; // @[Mux.scala 27:72]
  wire [63:0] _T_1735; // @[Mux.scala 27:72]
  wire [63:0] _GEN_503; // @[Mux.scala 27:72]
  wire [63:0] _T_1736; // @[Mux.scala 27:72]
  wire [63:0] _GEN_504; // @[Mux.scala 27:72]
  wire [63:0] _T_1737; // @[Mux.scala 27:72]
  wire [63:0] _T_1738; // @[Mux.scala 27:72]
  wire [63:0] _T_1739; // @[Mux.scala 27:72]
  wire [63:0] _GEN_505; // @[Mux.scala 27:72]
  wire [63:0] _T_1740; // @[Mux.scala 27:72]
  wire [63:0] _GEN_506; // @[Mux.scala 27:72]
  wire [63:0] _T_1741; // @[Mux.scala 27:72]
  wire [63:0] _GEN_507; // @[Mux.scala 27:72]
  wire [63:0] _T_1742; // @[Mux.scala 27:72]
  wire [63:0] _T_1743; // @[Mux.scala 27:72]
  wire [63:0] _T_1744; // @[Mux.scala 27:72]
  wire [63:0] _GEN_508; // @[Mux.scala 27:72]
  wire [63:0] _T_1832; // @[Mux.scala 27:72]
  wire [63:0] _T_1833; // @[Mux.scala 27:72]
  wire [63:0] _T_1834; // @[Mux.scala 27:72]
  wire [63:0] _T_1835; // @[Mux.scala 27:72]
  wire [63:0] _T_1836; // @[Mux.scala 27:72]
  wire [63:0] _T_1837; // @[Mux.scala 27:72]
  wire [63:0] _T_1838; // @[Mux.scala 27:72]
  wire [63:0] _T_1839; // @[Mux.scala 27:72]
  wire [63:0] _T_1840; // @[Mux.scala 27:72]
  wire [63:0] _T_1841; // @[Mux.scala 27:72]
  wire [63:0] _T_1842; // @[Mux.scala 27:72]
  wire [63:0] _T_1843; // @[Mux.scala 27:72]
  wire [63:0] _GEN_509; // @[Mux.scala 27:72]
  wire [63:0] _T_1844; // @[Mux.scala 27:72]
  wire [63:0] _T_1845; // @[Mux.scala 27:72]
  wire [63:0] _T_1846; // @[Mux.scala 27:72]
  wire [63:0] _T_1847; // @[Mux.scala 27:72]
  wire [63:0] _GEN_510; // @[Mux.scala 27:72]
  wire [63:0] _T_1849; // @[Mux.scala 27:72]
  wire [63:0] _GEN_511; // @[Mux.scala 27:72]
  wire [63:0] _T_1850; // @[Mux.scala 27:72]
  wire [63:0] _GEN_512; // @[Mux.scala 27:72]
  wire [63:0] _T_1851; // @[Mux.scala 27:72]
  wire [63:0] _GEN_513; // @[Mux.scala 27:72]
  wire [63:0] _T_1852; // @[Mux.scala 27:72]
  wire [63:0] _GEN_514; // @[Mux.scala 27:72]
  wire [63:0] _T_1853; // @[Mux.scala 27:72]
  wire [63:0] _GEN_515; // @[Mux.scala 27:72]
  wire [63:0] _T_1854; // @[Mux.scala 27:72]
  wire [63:0] _GEN_516; // @[Mux.scala 27:72]
  wire [63:0] _T_1855; // @[Mux.scala 27:72]
  wire [63:0] _GEN_517; // @[Mux.scala 27:72]
  wire [63:0] _T_1856; // @[Mux.scala 27:72]
  wire [63:0] _T_1865; // @[Mux.scala 27:72]
  wire [63:0] _T_1866; // @[Mux.scala 27:72]
  wire  _T_1872; // @[package.scala 15:47]
  wire  _T_1873; // @[package.scala 15:47]
  wire  _T_1874; // @[package.scala 15:47]
  wire [4:0] _T_3610; // @[CSR.scala 798:30]
  wire [4:0] _GEN_118; // @[CSR.scala 797:30]
  wire  _T_3614; // @[package.scala 64:59]
  wire  csr_wen; // @[package.scala 64:59]
  wire [102:0] _T_3628;
  wire  _T_3660; // @[CSR.scala 1073:35]
  wire  _T_3662; // @[CSR.scala 1094:73]
  wire [1:0] _GEN_124; // @[CSR.scala 812:39]
  wire  _T_3670; // @[CSR.scala 841:43]
  wire [3:0] _T_3673; // @[CSR.scala 843:38]
  wire [63:0] _GEN_518; // @[CSR.scala 843:32]
  wire [63:0] _T_3674; // @[CSR.scala 843:32]
  wire [63:0] _T_3676; // @[CSR.scala 843:55]
  wire [63:0] _T_3678; // @[CSR.scala 843:73]
  wire [63:0] _T_3679; // @[CSR.scala 843:62]
  wire [15:0] _T_3694; // @[CSR.scala 851:59]
  wire [15:0] _T_3696; // @[CSR.scala 1069:9]
  wire [63:0] _GEN_519; // @[CSR.scala 1069:34]
  wire [63:0] _T_3697; // @[CSR.scala 1069:34]
  wire [63:0] _T_3702; // @[CSR.scala 1069:43]
  wire [63:0] _T_3721; // @[CSR.scala 858:59]
  wire [63:0] _T_3723; // @[CSR.scala 1090:31]
  wire [63:0] _GEN_140; // @[CSR.scala 859:40]
  wire [63:0] _GEN_142; // @[CSR.scala 862:40]
  wire [63:0] _T_3725; // @[CSR.scala 863:62]
  wire [63:0] _GEN_145; // @[CSR.scala 1087:31]
  wire [63:0] _GEN_147; // @[CSR.scala 1087:31]
  wire [63:0] _GEN_150; // @[CSR.scala 876:40]
  wire [63:0] _GEN_152; // @[CSR.scala 877:40]
  wire [63:0] _GEN_154; // @[CSR.scala 878:38]
  wire [63:0] _GEN_155; // @[CSR.scala 878:38]
  wire  _T_3748; // @[CSR.scala 1073:35]
  wire [63:0] _GEN_161; // @[CSR.scala 893:42]
  wire [1:0] _GEN_165; // @[CSR.scala 897:41]
  wire [63:0] _T_3790; // @[CSR.scala 910:52]
  wire [63:0] _T_3791; // @[CSR.scala 910:78]
  wire [63:0] _T_3792; // @[CSR.scala 910:69]
  wire  _T_3816; // @[package.scala 15:47]
  wire  _T_3817; // @[package.scala 15:47]
  wire  _T_3818; // @[package.scala 64:59]
  wire [3:0] _T_3819; // @[CSR.scala 918:44]
  wire [63:0] _T_3822; // @[CSR.scala 924:64]
  wire [63:0] _T_3824; // @[CSR.scala 924:81]
  wire [63:0] _GEN_177; // @[CSR.scala 926:42]
  wire [63:0] _GEN_178; // @[CSR.scala 927:42]
  wire [63:0] _T_3828; // @[CSR.scala 928:64]
  wire [63:0] _GEN_183; // @[CSR.scala 932:44]
  wire [63:0] _GEN_184; // @[CSR.scala 935:44]
  wire  _T_3832; // @[CSR.scala 941:55]
  wire [63:0] _GEN_186; // @[CSR.scala 942:44]
  wire [63:0] _T_3866; // @[CSR.scala 1069:9]
  wire [63:0] _T_3867; // @[CSR.scala 1069:34]
  wire [63:0] _T_3872; // @[CSR.scala 1069:43]
  wire  _T_3890; // @[CSR.scala 951:38]
  wire  _GEN_187; // @[CSR.scala 953:51]
  wire [63:0] _GEN_203; // @[CSR.scala 941:70]
  wire  _T_3975; // @[CSR.scala 961:57]
  wire  _T_3985; // @[CSR.scala 965:31]
  wire  _T_3989; // @[PMP.scala 49:20]
  wire  _T_3990; // @[PMP.scala 51:62]
  wire  _T_3991; // @[PMP.scala 51:44]
  wire  _T_3993; // @[CSR.scala 970:45]
  wire [63:0] _GEN_258; // @[CSR.scala 970:71]
  wire  _T_3995; // @[CSR.scala 961:57]
  wire  _T_4005; // @[CSR.scala 965:31]
  wire  _T_4009; // @[PMP.scala 49:20]
  wire  _T_4010; // @[PMP.scala 51:62]
  wire  _T_4011; // @[PMP.scala 51:44]
  wire  _T_4013; // @[CSR.scala 970:45]
  wire [63:0] _GEN_265; // @[CSR.scala 970:71]
  wire  _T_4015; // @[CSR.scala 961:57]
  wire  _T_4025; // @[CSR.scala 965:31]
  wire  _T_4029; // @[PMP.scala 49:20]
  wire  _T_4030; // @[PMP.scala 51:62]
  wire  _T_4031; // @[PMP.scala 51:44]
  wire  _T_4033; // @[CSR.scala 970:45]
  wire [63:0] _GEN_272; // @[CSR.scala 970:71]
  wire  _T_4035; // @[CSR.scala 961:57]
  wire  _T_4045; // @[CSR.scala 965:31]
  wire  _T_4049; // @[PMP.scala 49:20]
  wire  _T_4050; // @[PMP.scala 51:62]
  wire  _T_4051; // @[PMP.scala 51:44]
  wire  _T_4053; // @[CSR.scala 970:45]
  wire [63:0] _GEN_279; // @[CSR.scala 970:71]
  wire  _T_4055; // @[CSR.scala 961:57]
  wire  _T_4065; // @[CSR.scala 965:31]
  wire  _T_4069; // @[PMP.scala 49:20]
  wire  _T_4070; // @[PMP.scala 51:62]
  wire  _T_4071; // @[PMP.scala 51:44]
  wire  _T_4073; // @[CSR.scala 970:45]
  wire [63:0] _GEN_286; // @[CSR.scala 970:71]
  wire  _T_4075; // @[CSR.scala 961:57]
  wire  _T_4085; // @[CSR.scala 965:31]
  wire  _T_4089; // @[PMP.scala 49:20]
  wire  _T_4090; // @[PMP.scala 51:62]
  wire  _T_4091; // @[PMP.scala 51:44]
  wire  _T_4093; // @[CSR.scala 970:45]
  wire [63:0] _GEN_293; // @[CSR.scala 970:71]
  wire  _T_4095; // @[CSR.scala 961:57]
  wire  _T_4105; // @[CSR.scala 965:31]
  wire  _T_4109; // @[PMP.scala 49:20]
  wire  _T_4110; // @[PMP.scala 51:62]
  wire  _T_4111; // @[PMP.scala 51:44]
  wire  _T_4113; // @[CSR.scala 970:45]
  wire [63:0] _GEN_300; // @[CSR.scala 970:71]
  wire  _T_4115; // @[CSR.scala 961:57]
  wire  _T_4125; // @[CSR.scala 965:31]
  wire  _T_4131; // @[PMP.scala 51:44]
  wire  _T_4133; // @[CSR.scala 970:45]
  wire [63:0] _GEN_307; // @[CSR.scala 970:71]
  wire [63:0] _T_4134; // @[CSR.scala 977:23]
  wire [63:0] _T_4136; // @[CSR.scala 977:38]
  wire [63:0] _T_4137; // @[CSR.scala 977:31]
  wire [1:0] _GEN_320; // @[CSR.scala 811:18]
  wire [63:0] _GEN_335; // @[CSR.scala 811:18]
  wire [63:0] _GEN_337; // @[CSR.scala 811:18]
  wire [63:0] _GEN_340; // @[CSR.scala 811:18]
  wire [63:0] _GEN_342; // @[CSR.scala 811:18]
  wire [63:0] _GEN_345; // @[CSR.scala 811:18]
  wire [63:0] _GEN_346; // @[CSR.scala 811:18]
  wire [63:0] _GEN_352; // @[CSR.scala 811:18]
  wire [63:0] _GEN_357; // @[CSR.scala 811:18]
  wire [63:0] _GEN_358; // @[CSR.scala 811:18]
  wire [63:0] _GEN_363; // @[CSR.scala 811:18]
  wire [63:0] _GEN_364; // @[CSR.scala 811:18]
  wire [63:0] _GEN_366; // @[CSR.scala 811:18]
  wire [63:0] _GEN_404; // @[CSR.scala 811:18]
  wire [63:0] _GEN_411; // @[CSR.scala 811:18]
  wire [63:0] _GEN_418; // @[CSR.scala 811:18]
  wire [63:0] _GEN_425; // @[CSR.scala 811:18]
  wire [63:0] _GEN_432; // @[CSR.scala 811:18]
  wire [63:0] _GEN_439; // @[CSR.scala 811:18]
  wire [63:0] _GEN_446; // @[CSR.scala 811:18]
  wire [63:0] _GEN_453; // @[CSR.scala 811:18]
  wire  _T_4163; // @[CSR.scala 1048:26]
  reg [19:0] CSRFile_state; // @[Register tracking CSRFile state]
  reg [31:0] _RAND_113;
  reg  CSRFile_cov [0:1048575]; // @[Coverage map for CSRFile]
  reg [31:0] _RAND_114;
  wire  CSRFile_cov_read_data; // @[Coverage map for CSRFile]
  wire [19:0] CSRFile_cov_read_addr; // @[Coverage map for CSRFile]
  wire  CSRFile_cov_write_data; // @[Coverage map for CSRFile]
  wire [19:0] CSRFile_cov_write_addr; // @[Coverage map for CSRFile]
  wire  CSRFile_cov_write_mask; // @[Coverage map for CSRFile]
  wire  CSRFile_cov_write_en; // @[Coverage map for CSRFile]
  reg [29:0] CSRFile_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_115;
  wire [1:0] reg_dcsr_ebreaku_shl;
  wire [19:0] reg_dcsr_ebreaku_pad;
  wire [2:0] reg_pmp_3_cfg_l_shl;
  wire [19:0] reg_pmp_3_cfg_l_pad;
  wire [7:0] reg_pmp_5_cfg_l_shl;
  wire [19:0] reg_pmp_5_cfg_l_pad;
  wire [13:0] reg_dcsr_ebreaks_shl;
  wire [19:0] reg_dcsr_ebreaks_pad;
  wire [14:0] reg_pmp_6_cfg_l_shl;
  wire [19:0] reg_pmp_6_cfg_l_pad;
  wire [10:0] reg_mip_ssip_shl;
  wire [19:0] reg_mip_ssip_pad;
  wire [6:0] reg_mip_seip_shl;
  wire [19:0] reg_mip_seip_pad;
  wire [7:0] reg_pmp_7_cfg_l_shl;
  wire [19:0] reg_pmp_7_cfg_l_pad;
  wire [19:0] reg_dcsr_ebreakm_shl;
  wire [19:0] reg_dcsr_ebreakm_pad;
  wire [4:0] reg_mstatus_spp_shl;
  wire [19:0] reg_mstatus_spp_pad;
  wire [14:0] reg_debug_shl;
  wire [19:0] reg_debug_pad;
  wire [19:0] reg_pmp_0_cfg_l_shl;
  wire [19:0] reg_pmp_0_cfg_l_pad;
  wire [12:0] reg_mstatus_mprv_shl;
  wire [19:0] reg_mstatus_mprv_pad;
  wire [19:0] reg_pmp_4_cfg_l_shl;
  wire [19:0] reg_pmp_4_cfg_l_pad;
  wire [19:0] reg_singleStepped_shl;
  wire [19:0] reg_singleStepped_pad;
  wire [4:0] reg_mstatus_mie_shl;
  wire [19:0] reg_mstatus_mie_pad;
  wire [19:0] reg_pmp_1_cfg_l_shl;
  wire [19:0] reg_pmp_1_cfg_l_pad;
  wire [8:0] reg_pmp_7_cfg_a_shl;
  wire [19:0] reg_pmp_7_cfg_a_pad;
  wire [1:0] reg_bp_0_control_dmode_shl;
  wire [19:0] reg_bp_0_control_dmode_pad;
  wire [11:0] reg_mip_stip_shl;
  wire [19:0] reg_mip_stip_pad;
  wire [15:0] reg_mstatus_sie_shl;
  wire [19:0] reg_mstatus_sie_pad;
  wire [5:0] reg_pmp_2_cfg_l_shl;
  wire [19:0] reg_pmp_2_cfg_l_pad;
  wire [3:0] reg_mstatus_prv_shl;
  wire [19:0] reg_mstatus_prv_pad;
  wire [19:0] CSRFile_xor7;
  wire [19:0] CSRFile_xor18;
  wire [19:0] CSRFile_xor8;
  wire [19:0] CSRFile_xor3;
  wire [19:0] CSRFile_xor20;
  wire [19:0] CSRFile_xor9;
  wire [19:0] CSRFile_xor22;
  wire [19:0] CSRFile_xor10;
  wire [19:0] CSRFile_xor4;
  wire [19:0] CSRFile_xor1;
  wire [19:0] CSRFile_xor24;
  wire [19:0] CSRFile_xor11;
  wire [19:0] CSRFile_xor26;
  wire [19:0] CSRFile_xor12;
  wire [19:0] CSRFile_xor5;
  wire [19:0] CSRFile_xor28;
  wire [19:0] CSRFile_xor13;
  wire [19:0] CSRFile_xor30;
  wire [19:0] CSRFile_xor14;
  wire [19:0] CSRFile_xor6;
  wire [19:0] CSRFile_xor2;
  wire [19:0] CSRFile_xor0;
  wire  stopEn0;
  wire  stopEn1;
  wire  CSRFile_or0;
  reg  CSRFile_metaAssert;
  reg [31:0] _RAND_116;
  assign system_insn = io_rw_cmd == 3'h4; // @[CSR.scala 589:31]
  assign _T_703 = {io_rw_addr, 20'h0}; // @[CSR.scala 601:28]
  assign _T_710 = _T_703 & 32'h12400000; // @[Decode.scala 14:65]
  assign _T_711 = _T_710 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_712 = _T_703 & 32'h40000000; // @[Decode.scala 14:65]
  assign _T_713 = _T_712 == 32'h40000000; // @[Decode.scala 14:121]
  assign _T_715 = _T_711 | _T_713; // @[Decode.scala 15:30]
  assign insn_ret = system_insn & _T_715; // @[CSR.scala 601:95]
  assign _GEN_93 = io_rw_addr[10] ? reg_dcsr_prv : reg_mstatus_mpp; // @[CSR.scala 745:53]
  assign _GEN_102 = io_rw_addr[9] ? _GEN_93 : {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 739:52]
  assign _T_704 = _T_703 & 32'h10100000; // @[Decode.scala 14:65]
  assign _T_705 = _T_704 == 32'h0; // @[Decode.scala 14:121]
  assign insn_call = system_insn & _T_705; // @[CSR.scala 601:95]
  assign _T_708 = _T_704 == 32'h100000; // @[Decode.scala 14:121]
  assign insn_break = system_insn & _T_708; // @[CSR.scala 601:95]
  assign _T_1197 = insn_call | insn_break; // @[CSR.scala 673:29]
  assign exception = _T_1197 | io_exception; // @[CSR.scala 673:43]
  assign _GEN_490 = {{2'd0}, reg_mstatus_prv}; // @[CSR.scala 637:36]
  assign _T_1143 = _GEN_490 + 4'h8; // @[CSR.scala 637:36]
  assign _T_1144 = insn_break ? 64'h3 : io_cause; // @[CSR.scala 638:14]
  assign cause = insn_call ? {{60'd0}, _T_1143} : _T_1144; // @[CSR.scala 637:8]
  assign cause_lsbs = cause[7:0]; // @[CSR.scala 639:25]
  assign _T_1146 = cause_lsbs == 8'he; // @[CSR.scala 640:53]
  assign causeIsDebugInt = cause[63] & _T_1146; // @[CSR.scala 640:39]
  assign _T_1158 = reg_singleStepped | causeIsDebugInt; // @[CSR.scala 643:60]
  assign causeIsDebugTrigger = ~cause[63] & _T_1146; // @[CSR.scala 641:44]
  assign _T_1159 = _T_1158 | causeIsDebugTrigger; // @[CSR.scala 643:79]
  assign _T_1152 = ~cause[63] & insn_break; // @[CSR.scala 642:42]
  assign _T_1155 = {reg_dcsr_ebreakm,1'h0,reg_dcsr_ebreaks,reg_dcsr_ebreaku}; // @[Cat.scala 29:58]
  assign _T_1156 = _T_1155 >> reg_mstatus_prv; // @[CSR.scala 642:134]
  assign causeIsDebugBreak = _T_1152 & _T_1156[0]; // @[CSR.scala 642:56]
  assign _T_1160 = _T_1159 | causeIsDebugBreak; // @[CSR.scala 643:102]
  assign trapToDebug = _T_1160 | reg_debug; // @[CSR.scala 643:123]
  assign _GEN_42 = reg_debug ? reg_mstatus_prv : 2'h3; // @[CSR.scala 690:25]
  assign _T_1163 = reg_mstatus_prv <= 2'h1; // @[CSR.scala 645:59]
  assign read_mideleg = reg_mideleg & 64'h222; // @[CSR.scala 373:36]
  assign _T_1166 = read_mideleg >> cause_lsbs; // @[CSR.scala 645:102]
  assign read_medeleg = reg_medeleg & 64'hb15d; // @[CSR.scala 377:36]
  assign _T_1168 = read_medeleg >> cause_lsbs; // @[CSR.scala 645:128]
  assign _T_1170 = cause[63] ? _T_1166[0] : _T_1168[0]; // @[CSR.scala 645:74]
  assign delegate = _T_1163 & _T_1170; // @[CSR.scala 645:68]
  assign _GEN_50 = delegate ? 2'h1 : 2'h3; // @[CSR.scala 697:27]
  assign _GEN_61 = trapToDebug ? _GEN_42 : _GEN_50; // @[CSR.scala 689:24]
  assign _GEN_79 = exception ? _GEN_61 : reg_mstatus_prv; // @[CSR.scala 688:20]
  assign new_prv = insn_ret ? _GEN_102 : _GEN_79; // @[CSR.scala 738:19]
  assign _T_1 = new_prv == 2'h2; // @[CSR.scala 1073:35]
  assign read_mcounteren = reg_mcounteren & 32'h7; // @[CSR.scala 393:30]
  assign read_scounteren = reg_scounteren & 32'h7; // @[CSR.scala 397:36]
  assign _GEN_491 = {{5'd0}, io_retire}; // @[Counters.scala 47:33]
  assign _T_40 = _T_39 + _GEN_491; // @[Counters.scala 47:33]
  assign _T_44 = _T_41 + 58'h1; // @[Counters.scala 52:43]
  assign _T_45 = {_T_41,_T_39}; // @[Cat.scala 29:58]
  assign _GEN_492 = {{5'd0}, ~io_csr_stall}; // @[Counters.scala 47:33]
  assign _T_48 = _T_47 + _GEN_492; // @[Counters.scala 47:33]
  assign _T_52 = _T_49 + 58'h1; // @[Counters.scala 52:43]
  assign _T_53 = {_T_49,_T_47}; // @[Cat.scala 29:58]
  assign mip_seip = reg_mip_seip | io_interrupts_seip; // @[CSR.scala 427:57]
  assign _T_61 = {io_interrupts_mtip,1'h0,reg_mip_stip,1'h0,io_interrupts_msip,1'h0,reg_mip_ssip,1'h0}; // @[CSR.scala 429:22]
  assign _T_69 = {4'h0,io_interrupts_meip,1'h0,mip_seip,1'h0,_T_61}; // @[CSR.scala 429:22]
  assign read_mip = _T_69 & 16'haaa; // @[CSR.scala 429:29]
  assign _GEN_493 = {{48'd0}, read_mip}; // @[CSR.scala 432:56]
  assign pending_interrupts = _GEN_493 & reg_mie; // @[CSR.scala 432:56]
  assign d_interrupts = {io_interrupts_debug, 14'h0}; // @[CSR.scala 433:42]
  assign _T_72 = _T_1163 | reg_mstatus_mie; // @[CSR.scala 434:51]
  assign _T_74 = ~pending_interrupts | read_mideleg; // @[CSR.scala 434:93]
  assign m_interrupts = _T_72 ? ~_T_74 : 64'h0; // @[CSR.scala 434:25]
  assign _T_76 = reg_mstatus_prv < 2'h1; // @[CSR.scala 435:42]
  assign _T_77 = reg_mstatus_prv == 2'h1; // @[CSR.scala 435:70]
  assign _T_78 = _T_77 & reg_mstatus_sie; // @[CSR.scala 435:80]
  assign _T_79 = _T_76 | _T_78; // @[CSR.scala 435:50]
  assign _T_80 = pending_interrupts & read_mideleg; // @[CSR.scala 435:120]
  assign s_interrupts = _T_79 ? _T_80 : 64'h0; // @[CSR.scala 435:25]
  assign _T_119 = d_interrupts[14] | d_interrupts[13]; // @[CSR.scala 1063:90]
  assign _T_120 = _T_119 | d_interrupts[12]; // @[CSR.scala 1063:90]
  assign _T_121 = _T_120 | d_interrupts[11]; // @[CSR.scala 1063:90]
  assign _T_122 = _T_121 | d_interrupts[3]; // @[CSR.scala 1063:90]
  assign _T_123 = _T_122 | d_interrupts[7]; // @[CSR.scala 1063:90]
  assign _T_124 = _T_123 | d_interrupts[9]; // @[CSR.scala 1063:90]
  assign _T_125 = _T_124 | d_interrupts[1]; // @[CSR.scala 1063:90]
  assign _T_126 = _T_125 | d_interrupts[5]; // @[CSR.scala 1063:90]
  assign _T_127 = _T_126 | d_interrupts[8]; // @[CSR.scala 1063:90]
  assign _T_128 = _T_127 | d_interrupts[0]; // @[CSR.scala 1063:90]
  assign _T_129 = _T_128 | d_interrupts[4]; // @[CSR.scala 1063:90]
  assign _T_130 = _T_129 | m_interrupts[15]; // @[CSR.scala 1063:90]
  assign _T_131 = _T_130 | m_interrupts[14]; // @[CSR.scala 1063:90]
  assign _T_132 = _T_131 | m_interrupts[13]; // @[CSR.scala 1063:90]
  assign _T_133 = _T_132 | m_interrupts[12]; // @[CSR.scala 1063:90]
  assign _T_134 = _T_133 | m_interrupts[11]; // @[CSR.scala 1063:90]
  assign _T_135 = _T_134 | m_interrupts[3]; // @[CSR.scala 1063:90]
  assign _T_136 = _T_135 | m_interrupts[7]; // @[CSR.scala 1063:90]
  assign _T_137 = _T_136 | m_interrupts[9]; // @[CSR.scala 1063:90]
  assign _T_138 = _T_137 | m_interrupts[1]; // @[CSR.scala 1063:90]
  assign _T_139 = _T_138 | m_interrupts[5]; // @[CSR.scala 1063:90]
  assign _T_140 = _T_139 | m_interrupts[8]; // @[CSR.scala 1063:90]
  assign _T_141 = _T_140 | m_interrupts[0]; // @[CSR.scala 1063:90]
  assign _T_142 = _T_141 | m_interrupts[4]; // @[CSR.scala 1063:90]
  assign _T_143 = _T_142 | s_interrupts[15]; // @[CSR.scala 1063:90]
  assign _T_144 = _T_143 | s_interrupts[14]; // @[CSR.scala 1063:90]
  assign _T_145 = _T_144 | s_interrupts[13]; // @[CSR.scala 1063:90]
  assign _T_146 = _T_145 | s_interrupts[12]; // @[CSR.scala 1063:90]
  assign _T_147 = _T_146 | s_interrupts[11]; // @[CSR.scala 1063:90]
  assign _T_148 = _T_147 | s_interrupts[3]; // @[CSR.scala 1063:90]
  assign _T_149 = _T_148 | s_interrupts[7]; // @[CSR.scala 1063:90]
  assign _T_150 = _T_149 | s_interrupts[9]; // @[CSR.scala 1063:90]
  assign _T_151 = _T_150 | s_interrupts[1]; // @[CSR.scala 1063:90]
  assign _T_152 = _T_151 | s_interrupts[5]; // @[CSR.scala 1063:90]
  assign _T_153 = _T_152 | s_interrupts[8]; // @[CSR.scala 1063:90]
  assign _T_154 = _T_153 | s_interrupts[0]; // @[CSR.scala 1063:90]
  assign anyInterrupt = _T_154 | s_interrupts[4]; // @[CSR.scala 1063:90]
  assign _T_193 = s_interrupts[0] ? 3'h0 : 3'h4; // @[Mux.scala 47:69]
  assign _T_194 = s_interrupts[8] ? 4'h8 : {{1'd0}, _T_193}; // @[Mux.scala 47:69]
  assign _T_195 = s_interrupts[5] ? 4'h5 : _T_194; // @[Mux.scala 47:69]
  assign _T_196 = s_interrupts[1] ? 4'h1 : _T_195; // @[Mux.scala 47:69]
  assign _T_197 = s_interrupts[9] ? 4'h9 : _T_196; // @[Mux.scala 47:69]
  assign _T_198 = s_interrupts[7] ? 4'h7 : _T_197; // @[Mux.scala 47:69]
  assign _T_199 = s_interrupts[3] ? 4'h3 : _T_198; // @[Mux.scala 47:69]
  assign _T_200 = s_interrupts[11] ? 4'hb : _T_199; // @[Mux.scala 47:69]
  assign _T_201 = s_interrupts[12] ? 4'hc : _T_200; // @[Mux.scala 47:69]
  assign _T_202 = s_interrupts[13] ? 4'hd : _T_201; // @[Mux.scala 47:69]
  assign _T_203 = s_interrupts[14] ? 4'he : _T_202; // @[Mux.scala 47:69]
  assign _T_204 = s_interrupts[15] ? 4'hf : _T_203; // @[Mux.scala 47:69]
  assign _T_205 = m_interrupts[4] ? 4'h4 : _T_204; // @[Mux.scala 47:69]
  assign _T_206 = m_interrupts[0] ? 4'h0 : _T_205; // @[Mux.scala 47:69]
  assign _T_207 = m_interrupts[8] ? 4'h8 : _T_206; // @[Mux.scala 47:69]
  assign _T_208 = m_interrupts[5] ? 4'h5 : _T_207; // @[Mux.scala 47:69]
  assign _T_209 = m_interrupts[1] ? 4'h1 : _T_208; // @[Mux.scala 47:69]
  assign _T_210 = m_interrupts[9] ? 4'h9 : _T_209; // @[Mux.scala 47:69]
  assign _T_211 = m_interrupts[7] ? 4'h7 : _T_210; // @[Mux.scala 47:69]
  assign _T_212 = m_interrupts[3] ? 4'h3 : _T_211; // @[Mux.scala 47:69]
  assign _T_213 = m_interrupts[11] ? 4'hb : _T_212; // @[Mux.scala 47:69]
  assign _T_214 = m_interrupts[12] ? 4'hc : _T_213; // @[Mux.scala 47:69]
  assign _T_215 = m_interrupts[13] ? 4'hd : _T_214; // @[Mux.scala 47:69]
  assign _T_216 = m_interrupts[14] ? 4'he : _T_215; // @[Mux.scala 47:69]
  assign _T_217 = m_interrupts[15] ? 4'hf : _T_216; // @[Mux.scala 47:69]
  assign _T_218 = d_interrupts[4] ? 4'h4 : _T_217; // @[Mux.scala 47:69]
  assign _T_219 = d_interrupts[0] ? 4'h0 : _T_218; // @[Mux.scala 47:69]
  assign _T_220 = d_interrupts[8] ? 4'h8 : _T_219; // @[Mux.scala 47:69]
  assign _T_221 = d_interrupts[5] ? 4'h5 : _T_220; // @[Mux.scala 47:69]
  assign _T_222 = d_interrupts[1] ? 4'h1 : _T_221; // @[Mux.scala 47:69]
  assign _T_223 = d_interrupts[9] ? 4'h9 : _T_222; // @[Mux.scala 47:69]
  assign _T_224 = d_interrupts[7] ? 4'h7 : _T_223; // @[Mux.scala 47:69]
  assign _T_225 = d_interrupts[3] ? 4'h3 : _T_224; // @[Mux.scala 47:69]
  assign _T_226 = d_interrupts[11] ? 4'hb : _T_225; // @[Mux.scala 47:69]
  assign _T_227 = d_interrupts[12] ? 4'hc : _T_226; // @[Mux.scala 47:69]
  assign _T_228 = d_interrupts[13] ? 4'hd : _T_227; // @[Mux.scala 47:69]
  assign whichInterrupt = d_interrupts[14] ? 4'he : _T_228; // @[Mux.scala 47:69]
  assign _GEN_494 = {{60'd0}, whichInterrupt}; // @[CSR.scala 438:43]
  assign _T_231 = anyInterrupt & ~io_singleStep; // @[CSR.scala 439:33]
  assign _T_232 = _T_231 | reg_singleStepped; // @[CSR.scala 439:51]
  assign _T_233 = reg_debug | io_status_cease; // @[CSR.scala 439:88]
  assign _T_238 = {reg_pmp_0_addr,reg_pmp_0_cfg_a[0]}; // @[Cat.scala 29:58]
  assign _T_241 = _T_238 + 31'h1; // @[PMP.scala 60:23]
  assign _T_243 = _T_238 & ~_T_241; // @[PMP.scala 60:14]
  assign _T_244 = {_T_243,2'h3}; // @[Cat.scala 29:58]
  assign _T_247 = {reg_pmp_1_addr,reg_pmp_1_cfg_a[0]}; // @[Cat.scala 29:58]
  assign _T_250 = _T_247 + 31'h1; // @[PMP.scala 60:23]
  assign _T_252 = _T_247 & ~_T_250; // @[PMP.scala 60:14]
  assign _T_253 = {_T_252,2'h3}; // @[Cat.scala 29:58]
  assign _T_256 = {reg_pmp_2_addr,reg_pmp_2_cfg_a[0]}; // @[Cat.scala 29:58]
  assign _T_259 = _T_256 + 31'h1; // @[PMP.scala 60:23]
  assign _T_261 = _T_256 & ~_T_259; // @[PMP.scala 60:14]
  assign _T_262 = {_T_261,2'h3}; // @[Cat.scala 29:58]
  assign _T_265 = {reg_pmp_3_addr,reg_pmp_3_cfg_a[0]}; // @[Cat.scala 29:58]
  assign _T_268 = _T_265 + 31'h1; // @[PMP.scala 60:23]
  assign _T_270 = _T_265 & ~_T_268; // @[PMP.scala 60:14]
  assign _T_271 = {_T_270,2'h3}; // @[Cat.scala 29:58]
  assign _T_274 = {reg_pmp_4_addr,reg_pmp_4_cfg_a[0]}; // @[Cat.scala 29:58]
  assign _T_277 = _T_274 + 31'h1; // @[PMP.scala 60:23]
  assign _T_279 = _T_274 & ~_T_277; // @[PMP.scala 60:14]
  assign _T_280 = {_T_279,2'h3}; // @[Cat.scala 29:58]
  assign _T_283 = {reg_pmp_5_addr,reg_pmp_5_cfg_a[0]}; // @[Cat.scala 29:58]
  assign _T_286 = _T_283 + 31'h1; // @[PMP.scala 60:23]
  assign _T_288 = _T_283 & ~_T_286; // @[PMP.scala 60:14]
  assign _T_289 = {_T_288,2'h3}; // @[Cat.scala 29:58]
  assign _T_292 = {reg_pmp_6_addr,reg_pmp_6_cfg_a[0]}; // @[Cat.scala 29:58]
  assign _T_295 = _T_292 + 31'h1; // @[PMP.scala 60:23]
  assign _T_297 = _T_292 & ~_T_295; // @[PMP.scala 60:14]
  assign _T_298 = {_T_297,2'h3}; // @[Cat.scala 29:58]
  assign _T_301 = {reg_pmp_7_addr,reg_pmp_7_cfg_a[0]}; // @[Cat.scala 29:58]
  assign _T_304 = _T_301 + 31'h1; // @[PMP.scala 60:23]
  assign _T_306 = _T_301 & ~_T_304; // @[PMP.scala 60:14]
  assign _T_307 = {_T_306,2'h3}; // @[Cat.scala 29:58]
  assign _T_313 = {io_status_hpie,io_status_spie,io_status_upie,io_status_mie,io_status_hie,io_status_sie,io_status_uie}; // @[CSR.scala 458:38]
  assign _T_321 = {io_status_sum,io_status_mprv,io_status_xs,io_status_fs,io_status_mpp,io_status_vs,io_status_spp,io_status_mpie,_T_313}; // @[CSR.scala 458:38]
  assign _T_328 = {io_status_sxl,io_status_uxl,io_status_sd_rv32,io_status_zero1,io_status_tsr,io_status_tw,io_status_tvm,io_status_mxr}; // @[CSR.scala 458:38]
  assign _T_337 = {io_status_debug,io_status_cease,io_status_wfi,io_status_isa,io_status_dprv,io_status_prv,io_status_sd,io_status_zero2,_T_328,_T_321}; // @[CSR.scala 458:38]
  assign read_mstatus = _T_337[63:0]; // @[CSR.scala 458:40]
  assign _T_339 = reg_mtvec[0] ? 8'hfe : 8'h2; // @[CSR.scala 1092:39]
  assign _T_341 = {{24'd0}, _T_339}; // @[package.scala 154:41]
  assign _T_343 = reg_mtvec & ~_T_341; // @[package.scala 154:35]
  assign read_mtvec = {32'h0,_T_343}; // @[Cat.scala 29:58]
  assign _T_345 = reg_stvec[0] ? 8'hfe : 8'h2; // @[CSR.scala 1092:39]
  assign _T_347 = {{31'd0}, _T_345}; // @[package.scala 154:41]
  assign _T_349 = reg_stvec & ~_T_347; // @[package.scala 154:35]
  assign _T_352 = _T_349[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  assign read_stvec = {_T_352,_T_349}; // @[Cat.scala 29:58]
  assign _T_358 = {reg_bp_0_control_m,1'h0,reg_bp_0_control_s,reg_bp_0_control_u,reg_bp_0_control_x,reg_bp_0_control_w,reg_bp_0_control_r}; // @[CSR.scala 464:48]
  assign _T_366 = {4'h2,reg_bp_0_control_dmode,46'h40000000000,reg_bp_0_control_action,1'h0,2'h0,reg_bp_0_control_tmatch,_T_358}; // @[CSR.scala 464:48]
  assign _T_369 = reg_bp_0_address[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  assign _T_370 = {_T_369,reg_bp_0_address}; // @[Cat.scala 29:58]
  assign _T_373 = reg_misa[2] ? 2'h1 : 2'h3; // @[CSR.scala 1091:36]
  assign _GEN_495 = {{38'd0}, _T_373}; // @[CSR.scala 1091:31]
  assign _T_374 = ~reg_mepc | _GEN_495; // @[CSR.scala 1091:31]
  assign _T_376 = ~_T_374[39]; // @[package.scala 112:38]
  assign _T_378 = _T_376 ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_379 = {_T_378,~_T_374}; // @[Cat.scala 29:58]
  assign _T_382 = reg_mtval[39] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_383 = {_T_382,reg_mtval}; // @[Cat.scala 29:58]
  assign _T_389 = {2'h0,1'h0,reg_dcsr_cause,3'h0,reg_dcsr_step,reg_dcsr_prv}; // @[CSR.scala 478:27]
  assign _T_396 = {4'h4,12'h0,reg_dcsr_ebreakm,1'h0,reg_dcsr_ebreaks,reg_dcsr_ebreaku,_T_389}; // @[CSR.scala 478:27]
  assign _T_400 = ~reg_dpc | _GEN_495; // @[CSR.scala 1091:31]
  assign _T_402 = ~_T_400[39]; // @[package.scala 112:38]
  assign _T_404 = _T_402 ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_405 = {_T_404,~_T_400}; // @[Cat.scala 29:58]
  assign read_fcsr = {reg_frm,reg_fflags}; // @[Cat.scala 29:58]
  assign _T_406 = reg_mie & read_mideleg; // @[CSR.scala 534:28]
  assign _T_407 = _GEN_493 & read_mideleg; // @[CSR.scala 535:29]
  assign _T_415 = {1'h0,io_status_spie,2'h0,1'h0,io_status_sie,1'h0}; // @[CSR.scala 549:57]
  assign _T_423 = {io_status_sum,1'h0,io_status_xs,io_status_fs,2'h0,io_status_vs,io_status_spp,1'h0,_T_415}; // @[CSR.scala 549:57]
  assign _T_430 = {2'h0,io_status_uxl,io_status_sd_rv32,8'h0,2'h0,1'h0,io_status_mxr}; // @[CSR.scala 549:57]
  assign _T_439 = {35'h0,4'h0,io_status_sd,27'h0,_T_430,_T_423}; // @[CSR.scala 549:57]
  assign _T_443 = reg_stval[39] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_444 = {_T_443,reg_stval}; // @[Cat.scala 29:58]
  assign _T_446 = {reg_satp_mode,16'h0,reg_satp_ppn}; // @[CSR.scala 555:43]
  assign _T_450 = ~reg_sepc | _GEN_495; // @[CSR.scala 1091:31]
  assign _T_452 = ~_T_450[39]; // @[package.scala 112:38]
  assign _T_454 = _T_452 ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_455 = {_T_454,~_T_450}; // @[Cat.scala 29:58]
  assign _T_461 = {reg_pmp_0_cfg_l,2'h0,reg_pmp_0_cfg_a,reg_pmp_0_cfg_x,reg_pmp_0_cfg_w,reg_pmp_0_cfg_r}; // @[package.scala 36:38]
  assign _T_471 = {reg_pmp_2_cfg_l,2'h0,reg_pmp_2_cfg_a,reg_pmp_2_cfg_x,reg_pmp_2_cfg_w,reg_pmp_2_cfg_r}; // @[package.scala 36:38]
  assign _T_481 = {reg_pmp_4_cfg_l,2'h0,reg_pmp_4_cfg_a,reg_pmp_4_cfg_x,reg_pmp_4_cfg_w,reg_pmp_4_cfg_r}; // @[package.scala 36:38]
  assign _T_491 = {reg_pmp_6_cfg_l,2'h0,reg_pmp_6_cfg_a,reg_pmp_6_cfg_x,reg_pmp_6_cfg_w,reg_pmp_6_cfg_r}; // @[package.scala 36:38]
  assign _T_497 = {reg_pmp_1_cfg_l,2'h0,reg_pmp_1_cfg_a,reg_pmp_1_cfg_x,reg_pmp_1_cfg_w,reg_pmp_1_cfg_r,_T_461}; // @[Cat.scala 29:58]
  assign _T_499 = {reg_pmp_3_cfg_l,2'h0,reg_pmp_3_cfg_a,reg_pmp_3_cfg_x,reg_pmp_3_cfg_w,reg_pmp_3_cfg_r,_T_471,_T_497}; // @[Cat.scala 29:58]
  assign _T_500 = {reg_pmp_5_cfg_l,2'h0,reg_pmp_5_cfg_a,reg_pmp_5_cfg_x,reg_pmp_5_cfg_w,reg_pmp_5_cfg_r,_T_481}; // @[Cat.scala 29:58]
  assign _T_503 = {reg_pmp_7_cfg_l,2'h0,reg_pmp_7_cfg_a,reg_pmp_7_cfg_x,reg_pmp_7_cfg_w,reg_pmp_7_cfg_r,_T_491,_T_500,_T_499}; // @[Cat.scala 29:58]
  assign _T_552 = io_rw_addr == 12'h7a1; // @[CSR.scala 586:73]
  assign _T_553 = io_rw_addr == 12'h7a2; // @[CSR.scala 586:73]
  assign _T_554 = io_rw_addr == 12'h301; // @[CSR.scala 586:73]
  assign _T_555 = io_rw_addr == 12'h300; // @[CSR.scala 586:73]
  assign _T_556 = io_rw_addr == 12'h305; // @[CSR.scala 586:73]
  assign _T_557 = io_rw_addr == 12'h344; // @[CSR.scala 586:73]
  assign _T_558 = io_rw_addr == 12'h304; // @[CSR.scala 586:73]
  assign _T_559 = io_rw_addr == 12'h340; // @[CSR.scala 586:73]
  assign _T_560 = io_rw_addr == 12'h341; // @[CSR.scala 586:73]
  assign _T_561 = io_rw_addr == 12'h343; // @[CSR.scala 586:73]
  assign _T_562 = io_rw_addr == 12'h342; // @[CSR.scala 586:73]
  assign _T_563 = io_rw_addr == 12'hf14; // @[CSR.scala 586:73]
  assign _T_564 = io_rw_addr == 12'h7b0; // @[CSR.scala 586:73]
  assign _T_565 = io_rw_addr == 12'h7b1; // @[CSR.scala 586:73]
  assign _T_566 = io_rw_addr == 12'h7b2; // @[CSR.scala 586:73]
  assign _T_567 = io_rw_addr == 12'h1; // @[CSR.scala 586:73]
  assign _T_568 = io_rw_addr == 12'h2; // @[CSR.scala 586:73]
  assign _T_569 = io_rw_addr == 12'h3; // @[CSR.scala 586:73]
  assign _T_570 = io_rw_addr == 12'hb00; // @[CSR.scala 586:73]
  assign _T_571 = io_rw_addr == 12'hb02; // @[CSR.scala 586:73]
  assign _T_659 = io_rw_addr == 12'h306; // @[CSR.scala 586:73]
  assign _T_660 = io_rw_addr == 12'hc00; // @[CSR.scala 586:73]
  assign _T_661 = io_rw_addr == 12'hc02; // @[CSR.scala 586:73]
  assign _T_662 = io_rw_addr == 12'h100; // @[CSR.scala 586:73]
  assign _T_663 = io_rw_addr == 12'h144; // @[CSR.scala 586:73]
  assign _T_664 = io_rw_addr == 12'h104; // @[CSR.scala 586:73]
  assign _T_665 = io_rw_addr == 12'h140; // @[CSR.scala 586:73]
  assign _T_666 = io_rw_addr == 12'h142; // @[CSR.scala 586:73]
  assign _T_667 = io_rw_addr == 12'h143; // @[CSR.scala 586:73]
  assign _T_668 = io_rw_addr == 12'h180; // @[CSR.scala 586:73]
  assign _T_669 = io_rw_addr == 12'h141; // @[CSR.scala 586:73]
  assign _T_670 = io_rw_addr == 12'h105; // @[CSR.scala 586:73]
  assign _T_671 = io_rw_addr == 12'h106; // @[CSR.scala 586:73]
  assign _T_672 = io_rw_addr == 12'h303; // @[CSR.scala 586:73]
  assign _T_673 = io_rw_addr == 12'h302; // @[CSR.scala 586:73]
  assign _T_674 = io_rw_addr == 12'h3a0; // @[CSR.scala 586:73]
  assign _T_676 = io_rw_addr == 12'h3b0; // @[CSR.scala 586:73]
  assign _T_677 = io_rw_addr == 12'h3b1; // @[CSR.scala 586:73]
  assign _T_678 = io_rw_addr == 12'h3b2; // @[CSR.scala 586:73]
  assign _T_679 = io_rw_addr == 12'h3b3; // @[CSR.scala 586:73]
  assign _T_680 = io_rw_addr == 12'h3b4; // @[CSR.scala 586:73]
  assign _T_681 = io_rw_addr == 12'h3b5; // @[CSR.scala 586:73]
  assign _T_682 = io_rw_addr == 12'h3b6; // @[CSR.scala 586:73]
  assign _T_683 = io_rw_addr == 12'h3b7; // @[CSR.scala 586:73]
  assign _T_692 = io_rw_addr == 12'h7c1; // @[CSR.scala 586:73]
  assign _T_693 = io_rw_addr == 12'hf12; // @[CSR.scala 586:73]
  assign _T_695 = io_rw_addr == 12'hf13; // @[CSR.scala 586:73]
  assign _T_697 = io_rw_cmd[1] ? io_rw_rdata : 64'h0; // @[CSR.scala 1069:9]
  assign _T_698 = _T_697 | io_rw_wdata; // @[CSR.scala 1069:34]
  assign _T_700 = &io_rw_cmd[1:0]; // @[CSR.scala 1069:59]
  assign _T_701 = _T_700 ? io_rw_wdata : 64'h0; // @[CSR.scala 1069:49]
  assign wdata = _T_698 & ~_T_701; // @[CSR.scala 1069:43]
  assign _T_716 = _T_703 & 32'h20200000; // @[Decode.scala 14:65]
  assign _T_717 = _T_716 == 32'h20000000; // @[Decode.scala 14:121]
  assign _T_719 = _T_703 & 32'h32200000; // @[Decode.scala 14:65]
  assign _T_720 = _T_719 == 32'h10000000; // @[Decode.scala 14:121]
  assign insn_cease = system_insn & _T_717; // @[CSR.scala 601:95]
  assign insn_wfi = system_insn & _T_720; // @[CSR.scala 601:95]
  assign _T_731 = {io_decode_0_csr, 20'h0}; // @[CSR.scala 608:30]
  assign _T_738 = _T_731 & 32'h12400000; // @[Decode.scala 14:65]
  assign _T_739 = _T_738 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_740 = _T_731 & 32'h40000000; // @[Decode.scala 14:65]
  assign _T_741 = _T_740 == 32'h40000000; // @[Decode.scala 14:121]
  assign _T_743 = _T_739 | _T_741; // @[Decode.scala 15:30]
  assign _T_747 = _T_731 & 32'h32200000; // @[Decode.scala 14:65]
  assign _T_748 = _T_747 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_750 = _T_731 & 32'h42000000; // @[Decode.scala 14:65]
  assign _T_751 = _T_750 == 32'h2000000; // @[Decode.scala 14:121]
  assign _T_759 = reg_mstatus_prv > 2'h1; // @[CSR.scala 610:63]
  assign _T_762 = _T_759 | ~reg_mstatus_tw; // @[CSR.scala 610:71]
  assign _T_766 = _T_759 | ~reg_mstatus_tvm; // @[CSR.scala 611:70]
  assign _T_770 = _T_759 | ~reg_mstatus_tsr; // @[CSR.scala 612:72]
  assign _T_773 = read_mcounteren >> io_decode_0_csr[4:0]; // @[CSR.scala 614:68]
  assign _T_775 = _T_759 | _T_773[0]; // @[CSR.scala 614:50]
  assign _T_776 = reg_mstatus_prv >= 2'h1; // @[CSR.scala 615:44]
  assign _T_778 = read_scounteren >> io_decode_0_csr[4:0]; // @[CSR.scala 615:71]
  assign _T_780 = _T_776 | _T_778[0]; // @[CSR.scala 615:53]
  assign _T_781 = _T_775 & _T_780; // @[CSR.scala 614:84]
  assign _T_782 = io_status_fs == 2'h0; // @[CSR.scala 616:39]
  assign _T_790 = io_decode_0_csr & 12'h900; // @[Decode.scala 14:65]
  assign _T_799 = reg_mstatus_prv < io_decode_0_csr[9:8]; // @[CSR.scala 620:44]
  assign _T_800 = io_decode_0_csr == 12'h7a0; // @[CSR.scala 604:99]
  assign _T_801 = io_decode_0_csr == 12'h7a1; // @[CSR.scala 604:99]
  assign _T_802 = io_decode_0_csr == 12'h7a2; // @[CSR.scala 604:99]
  assign _T_803 = io_decode_0_csr == 12'h301; // @[CSR.scala 604:99]
  assign _T_804 = io_decode_0_csr == 12'h300; // @[CSR.scala 604:99]
  assign _T_805 = io_decode_0_csr == 12'h305; // @[CSR.scala 604:99]
  assign _T_806 = io_decode_0_csr == 12'h344; // @[CSR.scala 604:99]
  assign _T_807 = io_decode_0_csr == 12'h304; // @[CSR.scala 604:99]
  assign _T_808 = io_decode_0_csr == 12'h340; // @[CSR.scala 604:99]
  assign _T_809 = io_decode_0_csr == 12'h341; // @[CSR.scala 604:99]
  assign _T_810 = io_decode_0_csr == 12'h343; // @[CSR.scala 604:99]
  assign _T_811 = io_decode_0_csr == 12'h342; // @[CSR.scala 604:99]
  assign _T_812 = io_decode_0_csr == 12'hf14; // @[CSR.scala 604:99]
  assign _T_813 = io_decode_0_csr == 12'h7b0; // @[CSR.scala 604:99]
  assign _T_814 = io_decode_0_csr == 12'h7b1; // @[CSR.scala 604:99]
  assign _T_815 = io_decode_0_csr == 12'h7b2; // @[CSR.scala 604:99]
  assign _T_816 = io_decode_0_csr == 12'h1; // @[CSR.scala 604:99]
  assign _T_817 = io_decode_0_csr == 12'h2; // @[CSR.scala 604:99]
  assign _T_818 = io_decode_0_csr == 12'h3; // @[CSR.scala 604:99]
  assign _T_819 = io_decode_0_csr == 12'hb00; // @[CSR.scala 604:99]
  assign _T_820 = io_decode_0_csr == 12'hb02; // @[CSR.scala 604:99]
  assign _T_821 = io_decode_0_csr == 12'h323; // @[CSR.scala 604:99]
  assign _T_822 = io_decode_0_csr == 12'hb03; // @[CSR.scala 604:99]
  assign _T_823 = io_decode_0_csr == 12'hc03; // @[CSR.scala 604:99]
  assign _T_824 = io_decode_0_csr == 12'h324; // @[CSR.scala 604:99]
  assign _T_825 = io_decode_0_csr == 12'hb04; // @[CSR.scala 604:99]
  assign _T_826 = io_decode_0_csr == 12'hc04; // @[CSR.scala 604:99]
  assign _T_827 = io_decode_0_csr == 12'h325; // @[CSR.scala 604:99]
  assign _T_828 = io_decode_0_csr == 12'hb05; // @[CSR.scala 604:99]
  assign _T_829 = io_decode_0_csr == 12'hc05; // @[CSR.scala 604:99]
  assign _T_830 = io_decode_0_csr == 12'h326; // @[CSR.scala 604:99]
  assign _T_831 = io_decode_0_csr == 12'hb06; // @[CSR.scala 604:99]
  assign _T_832 = io_decode_0_csr == 12'hc06; // @[CSR.scala 604:99]
  assign _T_833 = io_decode_0_csr == 12'h327; // @[CSR.scala 604:99]
  assign _T_834 = io_decode_0_csr == 12'hb07; // @[CSR.scala 604:99]
  assign _T_835 = io_decode_0_csr == 12'hc07; // @[CSR.scala 604:99]
  assign _T_836 = io_decode_0_csr == 12'h328; // @[CSR.scala 604:99]
  assign _T_837 = io_decode_0_csr == 12'hb08; // @[CSR.scala 604:99]
  assign _T_838 = io_decode_0_csr == 12'hc08; // @[CSR.scala 604:99]
  assign _T_839 = io_decode_0_csr == 12'h329; // @[CSR.scala 604:99]
  assign _T_840 = io_decode_0_csr == 12'hb09; // @[CSR.scala 604:99]
  assign _T_841 = io_decode_0_csr == 12'hc09; // @[CSR.scala 604:99]
  assign _T_842 = io_decode_0_csr == 12'h32a; // @[CSR.scala 604:99]
  assign _T_843 = io_decode_0_csr == 12'hb0a; // @[CSR.scala 604:99]
  assign _T_844 = io_decode_0_csr == 12'hc0a; // @[CSR.scala 604:99]
  assign _T_845 = io_decode_0_csr == 12'h32b; // @[CSR.scala 604:99]
  assign _T_846 = io_decode_0_csr == 12'hb0b; // @[CSR.scala 604:99]
  assign _T_847 = io_decode_0_csr == 12'hc0b; // @[CSR.scala 604:99]
  assign _T_848 = io_decode_0_csr == 12'h32c; // @[CSR.scala 604:99]
  assign _T_849 = io_decode_0_csr == 12'hb0c; // @[CSR.scala 604:99]
  assign _T_850 = io_decode_0_csr == 12'hc0c; // @[CSR.scala 604:99]
  assign _T_851 = io_decode_0_csr == 12'h32d; // @[CSR.scala 604:99]
  assign _T_852 = io_decode_0_csr == 12'hb0d; // @[CSR.scala 604:99]
  assign _T_853 = io_decode_0_csr == 12'hc0d; // @[CSR.scala 604:99]
  assign _T_854 = io_decode_0_csr == 12'h32e; // @[CSR.scala 604:99]
  assign _T_855 = io_decode_0_csr == 12'hb0e; // @[CSR.scala 604:99]
  assign _T_856 = io_decode_0_csr == 12'hc0e; // @[CSR.scala 604:99]
  assign _T_857 = io_decode_0_csr == 12'h32f; // @[CSR.scala 604:99]
  assign _T_858 = io_decode_0_csr == 12'hb0f; // @[CSR.scala 604:99]
  assign _T_859 = io_decode_0_csr == 12'hc0f; // @[CSR.scala 604:99]
  assign _T_860 = io_decode_0_csr == 12'h330; // @[CSR.scala 604:99]
  assign _T_861 = io_decode_0_csr == 12'hb10; // @[CSR.scala 604:99]
  assign _T_862 = io_decode_0_csr == 12'hc10; // @[CSR.scala 604:99]
  assign _T_863 = io_decode_0_csr == 12'h331; // @[CSR.scala 604:99]
  assign _T_864 = io_decode_0_csr == 12'hb11; // @[CSR.scala 604:99]
  assign _T_865 = io_decode_0_csr == 12'hc11; // @[CSR.scala 604:99]
  assign _T_866 = io_decode_0_csr == 12'h332; // @[CSR.scala 604:99]
  assign _T_867 = io_decode_0_csr == 12'hb12; // @[CSR.scala 604:99]
  assign _T_868 = io_decode_0_csr == 12'hc12; // @[CSR.scala 604:99]
  assign _T_869 = io_decode_0_csr == 12'h333; // @[CSR.scala 604:99]
  assign _T_870 = io_decode_0_csr == 12'hb13; // @[CSR.scala 604:99]
  assign _T_871 = io_decode_0_csr == 12'hc13; // @[CSR.scala 604:99]
  assign _T_872 = io_decode_0_csr == 12'h334; // @[CSR.scala 604:99]
  assign _T_873 = io_decode_0_csr == 12'hb14; // @[CSR.scala 604:99]
  assign _T_874 = io_decode_0_csr == 12'hc14; // @[CSR.scala 604:99]
  assign _T_875 = io_decode_0_csr == 12'h335; // @[CSR.scala 604:99]
  assign _T_876 = io_decode_0_csr == 12'hb15; // @[CSR.scala 604:99]
  assign _T_877 = io_decode_0_csr == 12'hc15; // @[CSR.scala 604:99]
  assign _T_878 = io_decode_0_csr == 12'h336; // @[CSR.scala 604:99]
  assign _T_879 = io_decode_0_csr == 12'hb16; // @[CSR.scala 604:99]
  assign _T_880 = io_decode_0_csr == 12'hc16; // @[CSR.scala 604:99]
  assign _T_881 = io_decode_0_csr == 12'h337; // @[CSR.scala 604:99]
  assign _T_882 = io_decode_0_csr == 12'hb17; // @[CSR.scala 604:99]
  assign _T_883 = io_decode_0_csr == 12'hc17; // @[CSR.scala 604:99]
  assign _T_884 = io_decode_0_csr == 12'h338; // @[CSR.scala 604:99]
  assign _T_885 = io_decode_0_csr == 12'hb18; // @[CSR.scala 604:99]
  assign _T_886 = io_decode_0_csr == 12'hc18; // @[CSR.scala 604:99]
  assign _T_887 = io_decode_0_csr == 12'h339; // @[CSR.scala 604:99]
  assign _T_888 = io_decode_0_csr == 12'hb19; // @[CSR.scala 604:99]
  assign _T_889 = io_decode_0_csr == 12'hc19; // @[CSR.scala 604:99]
  assign _T_890 = io_decode_0_csr == 12'h33a; // @[CSR.scala 604:99]
  assign _T_891 = io_decode_0_csr == 12'hb1a; // @[CSR.scala 604:99]
  assign _T_892 = io_decode_0_csr == 12'hc1a; // @[CSR.scala 604:99]
  assign _T_893 = io_decode_0_csr == 12'h33b; // @[CSR.scala 604:99]
  assign _T_894 = io_decode_0_csr == 12'hb1b; // @[CSR.scala 604:99]
  assign _T_895 = io_decode_0_csr == 12'hc1b; // @[CSR.scala 604:99]
  assign _T_896 = io_decode_0_csr == 12'h33c; // @[CSR.scala 604:99]
  assign _T_897 = io_decode_0_csr == 12'hb1c; // @[CSR.scala 604:99]
  assign _T_898 = io_decode_0_csr == 12'hc1c; // @[CSR.scala 604:99]
  assign _T_899 = io_decode_0_csr == 12'h33d; // @[CSR.scala 604:99]
  assign _T_900 = io_decode_0_csr == 12'hb1d; // @[CSR.scala 604:99]
  assign _T_901 = io_decode_0_csr == 12'hc1d; // @[CSR.scala 604:99]
  assign _T_902 = io_decode_0_csr == 12'h33e; // @[CSR.scala 604:99]
  assign _T_903 = io_decode_0_csr == 12'hb1e; // @[CSR.scala 604:99]
  assign _T_904 = io_decode_0_csr == 12'hc1e; // @[CSR.scala 604:99]
  assign _T_905 = io_decode_0_csr == 12'h33f; // @[CSR.scala 604:99]
  assign _T_906 = io_decode_0_csr == 12'hb1f; // @[CSR.scala 604:99]
  assign _T_907 = io_decode_0_csr == 12'hc1f; // @[CSR.scala 604:99]
  assign _T_908 = io_decode_0_csr == 12'h306; // @[CSR.scala 604:99]
  assign _T_909 = io_decode_0_csr == 12'hc00; // @[CSR.scala 604:99]
  assign _T_910 = io_decode_0_csr == 12'hc02; // @[CSR.scala 604:99]
  assign _T_911 = io_decode_0_csr == 12'h100; // @[CSR.scala 604:99]
  assign _T_912 = io_decode_0_csr == 12'h144; // @[CSR.scala 604:99]
  assign _T_913 = io_decode_0_csr == 12'h104; // @[CSR.scala 604:99]
  assign _T_914 = io_decode_0_csr == 12'h140; // @[CSR.scala 604:99]
  assign _T_915 = io_decode_0_csr == 12'h142; // @[CSR.scala 604:99]
  assign _T_916 = io_decode_0_csr == 12'h143; // @[CSR.scala 604:99]
  assign _T_917 = io_decode_0_csr == 12'h180; // @[CSR.scala 604:99]
  assign _T_918 = io_decode_0_csr == 12'h141; // @[CSR.scala 604:99]
  assign _T_919 = io_decode_0_csr == 12'h105; // @[CSR.scala 604:99]
  assign _T_920 = io_decode_0_csr == 12'h106; // @[CSR.scala 604:99]
  assign _T_921 = io_decode_0_csr == 12'h303; // @[CSR.scala 604:99]
  assign _T_922 = io_decode_0_csr == 12'h302; // @[CSR.scala 604:99]
  assign _T_923 = io_decode_0_csr == 12'h3a0; // @[CSR.scala 604:99]
  assign _T_924 = io_decode_0_csr == 12'h3a2; // @[CSR.scala 604:99]
  assign _T_925 = io_decode_0_csr == 12'h3b0; // @[CSR.scala 604:99]
  assign _T_926 = io_decode_0_csr == 12'h3b1; // @[CSR.scala 604:99]
  assign _T_927 = io_decode_0_csr == 12'h3b2; // @[CSR.scala 604:99]
  assign _T_928 = io_decode_0_csr == 12'h3b3; // @[CSR.scala 604:99]
  assign _T_929 = io_decode_0_csr == 12'h3b4; // @[CSR.scala 604:99]
  assign _T_930 = io_decode_0_csr == 12'h3b5; // @[CSR.scala 604:99]
  assign _T_931 = io_decode_0_csr == 12'h3b6; // @[CSR.scala 604:99]
  assign _T_932 = io_decode_0_csr == 12'h3b7; // @[CSR.scala 604:99]
  assign _T_933 = io_decode_0_csr == 12'h3b8; // @[CSR.scala 604:99]
  assign _T_934 = io_decode_0_csr == 12'h3b9; // @[CSR.scala 604:99]
  assign _T_935 = io_decode_0_csr == 12'h3ba; // @[CSR.scala 604:99]
  assign _T_936 = io_decode_0_csr == 12'h3bb; // @[CSR.scala 604:99]
  assign _T_937 = io_decode_0_csr == 12'h3bc; // @[CSR.scala 604:99]
  assign _T_938 = io_decode_0_csr == 12'h3bd; // @[CSR.scala 604:99]
  assign _T_939 = io_decode_0_csr == 12'h3be; // @[CSR.scala 604:99]
  assign _T_940 = io_decode_0_csr == 12'h3bf; // @[CSR.scala 604:99]
  assign _T_941 = io_decode_0_csr == 12'h7c1; // @[CSR.scala 604:99]
  assign _T_942 = io_decode_0_csr == 12'hf12; // @[CSR.scala 604:99]
  assign _T_943 = io_decode_0_csr == 12'hf11; // @[CSR.scala 604:99]
  assign _T_944 = io_decode_0_csr == 12'hf13; // @[CSR.scala 604:99]
  assign _T_945 = _T_800 | _T_801; // @[CSR.scala 604:115]
  assign _T_946 = _T_945 | _T_802; // @[CSR.scala 604:115]
  assign _T_947 = _T_946 | _T_803; // @[CSR.scala 604:115]
  assign _T_948 = _T_947 | _T_804; // @[CSR.scala 604:115]
  assign _T_949 = _T_948 | _T_805; // @[CSR.scala 604:115]
  assign _T_950 = _T_949 | _T_806; // @[CSR.scala 604:115]
  assign _T_951 = _T_950 | _T_807; // @[CSR.scala 604:115]
  assign _T_952 = _T_951 | _T_808; // @[CSR.scala 604:115]
  assign _T_953 = _T_952 | _T_809; // @[CSR.scala 604:115]
  assign _T_954 = _T_953 | _T_810; // @[CSR.scala 604:115]
  assign _T_955 = _T_954 | _T_811; // @[CSR.scala 604:115]
  assign _T_956 = _T_955 | _T_812; // @[CSR.scala 604:115]
  assign _T_957 = _T_956 | _T_813; // @[CSR.scala 604:115]
  assign _T_958 = _T_957 | _T_814; // @[CSR.scala 604:115]
  assign _T_959 = _T_958 | _T_815; // @[CSR.scala 604:115]
  assign _T_960 = _T_959 | _T_816; // @[CSR.scala 604:115]
  assign _T_961 = _T_960 | _T_817; // @[CSR.scala 604:115]
  assign _T_962 = _T_961 | _T_818; // @[CSR.scala 604:115]
  assign _T_963 = _T_962 | _T_819; // @[CSR.scala 604:115]
  assign _T_964 = _T_963 | _T_820; // @[CSR.scala 604:115]
  assign _T_965 = _T_964 | _T_821; // @[CSR.scala 604:115]
  assign _T_966 = _T_965 | _T_822; // @[CSR.scala 604:115]
  assign _T_967 = _T_966 | _T_823; // @[CSR.scala 604:115]
  assign _T_968 = _T_967 | _T_824; // @[CSR.scala 604:115]
  assign _T_969 = _T_968 | _T_825; // @[CSR.scala 604:115]
  assign _T_970 = _T_969 | _T_826; // @[CSR.scala 604:115]
  assign _T_971 = _T_970 | _T_827; // @[CSR.scala 604:115]
  assign _T_972 = _T_971 | _T_828; // @[CSR.scala 604:115]
  assign _T_973 = _T_972 | _T_829; // @[CSR.scala 604:115]
  assign _T_974 = _T_973 | _T_830; // @[CSR.scala 604:115]
  assign _T_975 = _T_974 | _T_831; // @[CSR.scala 604:115]
  assign _T_976 = _T_975 | _T_832; // @[CSR.scala 604:115]
  assign _T_977 = _T_976 | _T_833; // @[CSR.scala 604:115]
  assign _T_978 = _T_977 | _T_834; // @[CSR.scala 604:115]
  assign _T_979 = _T_978 | _T_835; // @[CSR.scala 604:115]
  assign _T_980 = _T_979 | _T_836; // @[CSR.scala 604:115]
  assign _T_981 = _T_980 | _T_837; // @[CSR.scala 604:115]
  assign _T_982 = _T_981 | _T_838; // @[CSR.scala 604:115]
  assign _T_983 = _T_982 | _T_839; // @[CSR.scala 604:115]
  assign _T_984 = _T_983 | _T_840; // @[CSR.scala 604:115]
  assign _T_985 = _T_984 | _T_841; // @[CSR.scala 604:115]
  assign _T_986 = _T_985 | _T_842; // @[CSR.scala 604:115]
  assign _T_987 = _T_986 | _T_843; // @[CSR.scala 604:115]
  assign _T_988 = _T_987 | _T_844; // @[CSR.scala 604:115]
  assign _T_989 = _T_988 | _T_845; // @[CSR.scala 604:115]
  assign _T_990 = _T_989 | _T_846; // @[CSR.scala 604:115]
  assign _T_991 = _T_990 | _T_847; // @[CSR.scala 604:115]
  assign _T_992 = _T_991 | _T_848; // @[CSR.scala 604:115]
  assign _T_993 = _T_992 | _T_849; // @[CSR.scala 604:115]
  assign _T_994 = _T_993 | _T_850; // @[CSR.scala 604:115]
  assign _T_995 = _T_994 | _T_851; // @[CSR.scala 604:115]
  assign _T_996 = _T_995 | _T_852; // @[CSR.scala 604:115]
  assign _T_997 = _T_996 | _T_853; // @[CSR.scala 604:115]
  assign _T_998 = _T_997 | _T_854; // @[CSR.scala 604:115]
  assign _T_999 = _T_998 | _T_855; // @[CSR.scala 604:115]
  assign _T_1000 = _T_999 | _T_856; // @[CSR.scala 604:115]
  assign _T_1001 = _T_1000 | _T_857; // @[CSR.scala 604:115]
  assign _T_1002 = _T_1001 | _T_858; // @[CSR.scala 604:115]
  assign _T_1003 = _T_1002 | _T_859; // @[CSR.scala 604:115]
  assign _T_1004 = _T_1003 | _T_860; // @[CSR.scala 604:115]
  assign _T_1005 = _T_1004 | _T_861; // @[CSR.scala 604:115]
  assign _T_1006 = _T_1005 | _T_862; // @[CSR.scala 604:115]
  assign _T_1007 = _T_1006 | _T_863; // @[CSR.scala 604:115]
  assign _T_1008 = _T_1007 | _T_864; // @[CSR.scala 604:115]
  assign _T_1009 = _T_1008 | _T_865; // @[CSR.scala 604:115]
  assign _T_1010 = _T_1009 | _T_866; // @[CSR.scala 604:115]
  assign _T_1011 = _T_1010 | _T_867; // @[CSR.scala 604:115]
  assign _T_1012 = _T_1011 | _T_868; // @[CSR.scala 604:115]
  assign _T_1013 = _T_1012 | _T_869; // @[CSR.scala 604:115]
  assign _T_1014 = _T_1013 | _T_870; // @[CSR.scala 604:115]
  assign _T_1015 = _T_1014 | _T_871; // @[CSR.scala 604:115]
  assign _T_1016 = _T_1015 | _T_872; // @[CSR.scala 604:115]
  assign _T_1017 = _T_1016 | _T_873; // @[CSR.scala 604:115]
  assign _T_1018 = _T_1017 | _T_874; // @[CSR.scala 604:115]
  assign _T_1019 = _T_1018 | _T_875; // @[CSR.scala 604:115]
  assign _T_1020 = _T_1019 | _T_876; // @[CSR.scala 604:115]
  assign _T_1021 = _T_1020 | _T_877; // @[CSR.scala 604:115]
  assign _T_1022 = _T_1021 | _T_878; // @[CSR.scala 604:115]
  assign _T_1023 = _T_1022 | _T_879; // @[CSR.scala 604:115]
  assign _T_1024 = _T_1023 | _T_880; // @[CSR.scala 604:115]
  assign _T_1025 = _T_1024 | _T_881; // @[CSR.scala 604:115]
  assign _T_1026 = _T_1025 | _T_882; // @[CSR.scala 604:115]
  assign _T_1027 = _T_1026 | _T_883; // @[CSR.scala 604:115]
  assign _T_1028 = _T_1027 | _T_884; // @[CSR.scala 604:115]
  assign _T_1029 = _T_1028 | _T_885; // @[CSR.scala 604:115]
  assign _T_1030 = _T_1029 | _T_886; // @[CSR.scala 604:115]
  assign _T_1031 = _T_1030 | _T_887; // @[CSR.scala 604:115]
  assign _T_1032 = _T_1031 | _T_888; // @[CSR.scala 604:115]
  assign _T_1033 = _T_1032 | _T_889; // @[CSR.scala 604:115]
  assign _T_1034 = _T_1033 | _T_890; // @[CSR.scala 604:115]
  assign _T_1035 = _T_1034 | _T_891; // @[CSR.scala 604:115]
  assign _T_1036 = _T_1035 | _T_892; // @[CSR.scala 604:115]
  assign _T_1037 = _T_1036 | _T_893; // @[CSR.scala 604:115]
  assign _T_1038 = _T_1037 | _T_894; // @[CSR.scala 604:115]
  assign _T_1039 = _T_1038 | _T_895; // @[CSR.scala 604:115]
  assign _T_1040 = _T_1039 | _T_896; // @[CSR.scala 604:115]
  assign _T_1041 = _T_1040 | _T_897; // @[CSR.scala 604:115]
  assign _T_1042 = _T_1041 | _T_898; // @[CSR.scala 604:115]
  assign _T_1043 = _T_1042 | _T_899; // @[CSR.scala 604:115]
  assign _T_1044 = _T_1043 | _T_900; // @[CSR.scala 604:115]
  assign _T_1045 = _T_1044 | _T_901; // @[CSR.scala 604:115]
  assign _T_1046 = _T_1045 | _T_902; // @[CSR.scala 604:115]
  assign _T_1047 = _T_1046 | _T_903; // @[CSR.scala 604:115]
  assign _T_1048 = _T_1047 | _T_904; // @[CSR.scala 604:115]
  assign _T_1049 = _T_1048 | _T_905; // @[CSR.scala 604:115]
  assign _T_1050 = _T_1049 | _T_906; // @[CSR.scala 604:115]
  assign _T_1051 = _T_1050 | _T_907; // @[CSR.scala 604:115]
  assign _T_1052 = _T_1051 | _T_908; // @[CSR.scala 604:115]
  assign _T_1053 = _T_1052 | _T_909; // @[CSR.scala 604:115]
  assign _T_1054 = _T_1053 | _T_910; // @[CSR.scala 604:115]
  assign _T_1055 = _T_1054 | _T_911; // @[CSR.scala 604:115]
  assign _T_1056 = _T_1055 | _T_912; // @[CSR.scala 604:115]
  assign _T_1057 = _T_1056 | _T_913; // @[CSR.scala 604:115]
  assign _T_1058 = _T_1057 | _T_914; // @[CSR.scala 604:115]
  assign _T_1059 = _T_1058 | _T_915; // @[CSR.scala 604:115]
  assign _T_1060 = _T_1059 | _T_916; // @[CSR.scala 604:115]
  assign _T_1061 = _T_1060 | _T_917; // @[CSR.scala 604:115]
  assign _T_1062 = _T_1061 | _T_918; // @[CSR.scala 604:115]
  assign _T_1063 = _T_1062 | _T_919; // @[CSR.scala 604:115]
  assign _T_1064 = _T_1063 | _T_920; // @[CSR.scala 604:115]
  assign _T_1065 = _T_1064 | _T_921; // @[CSR.scala 604:115]
  assign _T_1066 = _T_1065 | _T_922; // @[CSR.scala 604:115]
  assign _T_1067 = _T_1066 | _T_923; // @[CSR.scala 604:115]
  assign _T_1068 = _T_1067 | _T_924; // @[CSR.scala 604:115]
  assign _T_1069 = _T_1068 | _T_925; // @[CSR.scala 604:115]
  assign _T_1070 = _T_1069 | _T_926; // @[CSR.scala 604:115]
  assign _T_1071 = _T_1070 | _T_927; // @[CSR.scala 604:115]
  assign _T_1072 = _T_1071 | _T_928; // @[CSR.scala 604:115]
  assign _T_1073 = _T_1072 | _T_929; // @[CSR.scala 604:115]
  assign _T_1074 = _T_1073 | _T_930; // @[CSR.scala 604:115]
  assign _T_1075 = _T_1074 | _T_931; // @[CSR.scala 604:115]
  assign _T_1076 = _T_1075 | _T_932; // @[CSR.scala 604:115]
  assign _T_1077 = _T_1076 | _T_933; // @[CSR.scala 604:115]
  assign _T_1078 = _T_1077 | _T_934; // @[CSR.scala 604:115]
  assign _T_1079 = _T_1078 | _T_935; // @[CSR.scala 604:115]
  assign _T_1080 = _T_1079 | _T_936; // @[CSR.scala 604:115]
  assign _T_1081 = _T_1080 | _T_937; // @[CSR.scala 604:115]
  assign _T_1082 = _T_1081 | _T_938; // @[CSR.scala 604:115]
  assign _T_1083 = _T_1082 | _T_939; // @[CSR.scala 604:115]
  assign _T_1084 = _T_1083 | _T_940; // @[CSR.scala 604:115]
  assign _T_1085 = _T_1084 | _T_941; // @[CSR.scala 604:115]
  assign _T_1086 = _T_1085 | _T_942; // @[CSR.scala 604:115]
  assign _T_1087 = _T_1086 | _T_943; // @[CSR.scala 604:115]
  assign _T_1088 = _T_1087 | _T_944; // @[CSR.scala 604:115]
  assign _T_1090 = _T_799 | ~_T_1088; // @[CSR.scala 620:62]
  assign _T_1093 = _T_917 & ~_T_766; // @[CSR.scala 622:32]
  assign _T_1094 = _T_1090 | _T_1093; // @[CSR.scala 621:32]
  assign _T_1095 = io_decode_0_csr >= 12'hc00; // @[package.scala 185:47]
  assign _T_1096 = io_decode_0_csr < 12'hc20; // @[package.scala 185:60]
  assign _T_1097 = _T_1095 & _T_1096; // @[package.scala 185:55]
  assign _T_1098 = io_decode_0_csr >= 12'hc80; // @[package.scala 185:47]
  assign _T_1099 = io_decode_0_csr < 12'hca0; // @[package.scala 185:60]
  assign _T_1100 = _T_1098 & _T_1099; // @[package.scala 185:55]
  assign _T_1101 = _T_1097 | _T_1100; // @[CSR.scala 623:66]
  assign _T_1103 = _T_1101 & ~_T_781; // @[CSR.scala 623:130]
  assign _T_1104 = _T_1094 | _T_1103; // @[CSR.scala 622:53]
  assign _T_1105 = io_decode_0_csr & 12'hc10; // @[Decode.scala 14:65]
  assign _T_1106 = _T_1105 == 12'h410; // @[Decode.scala 14:121]
  assign _T_1110 = _T_1106 & ~reg_debug; // @[CSR.scala 624:42]
  assign _T_1111 = _T_1104 | _T_1110; // @[CSR.scala 623:148]
  assign _T_1114 = io_decode_0_fp_csr & io_decode_0_fp_illegal; // @[CSR.scala 626:21]
  assign _T_1118 = io_decode_0_csr >= 12'h340; // @[CSR.scala 628:40]
  assign _T_1119 = io_decode_0_csr <= 12'h343; // @[CSR.scala 628:71]
  assign _T_1120 = _T_1118 & _T_1119; // @[CSR.scala 628:57]
  assign _T_1121 = io_decode_0_csr >= 12'h140; // @[CSR.scala 628:99]
  assign _T_1122 = io_decode_0_csr <= 12'h143; // @[CSR.scala 628:130]
  assign _T_1123 = _T_1121 & _T_1122; // @[CSR.scala 628:116]
  assign _T_1124 = _T_1120 | _T_1123; // @[CSR.scala 628:85]
  assign _T_1129 = _T_748 & ~_T_762; // @[CSR.scala 630:14]
  assign _T_1130 = _T_799 | _T_1129; // @[CSR.scala 629:64]
  assign _T_1132 = _T_743 & ~_T_770; // @[CSR.scala 631:14]
  assign _T_1133 = _T_1130 | _T_1132; // @[CSR.scala 630:28]
  assign _T_1135 = _T_743 & io_decode_0_csr[10]; // @[CSR.scala 632:14]
  assign _T_1137 = _T_1135 & ~reg_debug; // @[CSR.scala 632:32]
  assign _T_1138 = _T_1133 | _T_1137; // @[CSR.scala 631:29]
  assign _T_1140 = _T_751 & ~_T_766; // @[CSR.scala 633:17]
  assign _T_1162 = insn_break ? 12'h800 : 12'h808; // @[CSR.scala 644:37]
  assign debugTVec = reg_debug ? _T_1162 : 12'h800; // @[CSR.scala 644:22]
  assign _T_1171 = delegate ? read_stvec : read_mtvec; // @[CSR.scala 652:19]
  assign _T_1173 = {cause[5:0], 2'h0}; // @[CSR.scala 653:59]
  assign _T_1175 = {_T_1171[63:8],_T_1173}; // @[Cat.scala 29:58]
  assign _T_1178 = _T_1171[0] & cause[63]; // @[CSR.scala 655:28]
  assign _T_1180 = cause_lsbs[7:6] == 2'h0; // @[CSR.scala 655:94]
  assign _T_1181 = _T_1178 & _T_1180; // @[CSR.scala 655:55]
  assign _T_1183 = {_T_1171[63:2], 2'h0}; // @[CSR.scala 656:56]
  assign notDebugTVec = _T_1181 ? _T_1175 : _T_1183; // @[CSR.scala 656:8]
  assign tvec = trapToDebug ? {{52'd0}, debugTVec} : notDebugTVec; // @[CSR.scala 658:17]
  assign _T_1188 = &io_status_fs; // @[CSR.scala 664:32]
  assign _T_1189 = &io_status_xs; // @[CSR.scala 664:53]
  assign _T_1190 = _T_1188 | _T_1189; // @[CSR.scala 664:37]
  assign _T_1191 = &io_status_vs; // @[CSR.scala 664:74]
  assign _T_1194 = reg_mstatus_mprv & ~reg_debug; // @[CSR.scala 669:53]
  assign _T_1198 = insn_ret + insn_call; // @[Bitwise.scala 47:55]
  assign _T_1200 = insn_break + io_exception; // @[Bitwise.scala 47:55]
  assign _T_1202 = _T_1198 + _T_1200; // @[Bitwise.scala 47:55]
  assign _T_1204 = _T_1202 <= 3'h1; // @[CSR.scala 674:79]
  assign _T_1206 = _T_1204 | reset; // @[CSR.scala 674:9]
  assign _T_1209 = insn_wfi & ~io_singleStep; // @[CSR.scala 676:18]
  assign _T_1211 = _T_1209 & ~reg_debug; // @[CSR.scala 676:36]
  assign _GEN_34 = _T_1211 | reg_wfi; // @[CSR.scala 676:51]
  assign _T_1212 = |pending_interrupts; // @[CSR.scala 677:28]
  assign _T_1213 = _T_1212 | io_interrupts_debug; // @[CSR.scala 677:32]
  assign _T_1214 = _T_1213 | exception; // @[CSR.scala 677:55]
  assign _T_1216 = io_retire | exception; // @[CSR.scala 679:22]
  assign _GEN_36 = _T_1216 | reg_singleStepped; // @[CSR.scala 679:36]
  assign _T_1226 = ~reg_singleStepped | ~io_retire; // @[CSR.scala 682:29]
  assign _T_1228 = _T_1226 | reset; // @[CSR.scala 682:9]
  assign _T_1231 = ~io_pc | 40'h1; // @[CSR.scala 1090:31]
  assign epc = ~_T_1231; // @[CSR.scala 1090:26]
  assign _T_1233 = causeIsDebugTrigger ? 2'h2 : 2'h1; // @[CSR.scala 693:86]
  assign _T_1234 = causeIsDebugInt ? 2'h3 : _T_1233; // @[CSR.scala 693:56]
  assign _GEN_38 = ~reg_debug | reg_debug; // @[CSR.scala 690:25]
  assign _GEN_39 = reg_debug ? reg_dpc : epc; // @[CSR.scala 690:25]
  assign _GEN_43 = delegate ? epc : reg_sepc; // @[CSR.scala 697:27]
  assign _GEN_47 = delegate ? reg_mstatus_sie : reg_mstatus_spie; // @[CSR.scala 697:27]
  assign _GEN_48 = delegate ? reg_mstatus_prv : {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 697:27]
  assign _GEN_51 = delegate ? reg_mepc : epc; // @[CSR.scala 697:27]
  assign _GEN_54 = delegate ? reg_mstatus_mpie : reg_mstatus_mie; // @[CSR.scala 697:27]
  assign _GEN_55 = delegate ? reg_mstatus_mpp : reg_mstatus_prv; // @[CSR.scala 697:27]
  assign _GEN_56 = delegate & reg_mstatus_mie; // @[CSR.scala 697:27]
  assign _GEN_58 = trapToDebug ? _GEN_39 : reg_dpc; // @[CSR.scala 689:24]
  assign _GEN_62 = trapToDebug ? reg_sepc : _GEN_43; // @[CSR.scala 689:24]
  assign _GEN_66 = trapToDebug ? reg_mstatus_spie : _GEN_47; // @[CSR.scala 689:24]
  assign _GEN_67 = trapToDebug ? {{1'd0}, reg_mstatus_spp} : _GEN_48; // @[CSR.scala 689:24]
  assign _GEN_69 = trapToDebug ? reg_mepc : _GEN_51; // @[CSR.scala 689:24]
  assign _GEN_72 = trapToDebug ? reg_mstatus_mpie : _GEN_54; // @[CSR.scala 689:24]
  assign _GEN_73 = trapToDebug ? reg_mstatus_mpp : _GEN_55; // @[CSR.scala 689:24]
  assign _GEN_74 = trapToDebug ? reg_mstatus_mie : _GEN_56; // @[CSR.scala 689:24]
  assign _GEN_76 = exception ? _GEN_58 : reg_dpc; // @[CSR.scala 688:20]
  assign _GEN_80 = exception ? _GEN_62 : reg_sepc; // @[CSR.scala 688:20]
  assign _GEN_84 = exception ? _GEN_66 : reg_mstatus_spie; // @[CSR.scala 688:20]
  assign _GEN_85 = exception ? _GEN_67 : {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 688:20]
  assign _GEN_87 = exception ? _GEN_69 : reg_mepc; // @[CSR.scala 688:20]
  assign _GEN_90 = exception ? _GEN_72 : reg_mstatus_mpie; // @[CSR.scala 688:20]
  assign _GEN_91 = exception ? _GEN_73 : reg_mstatus_mpp; // @[CSR.scala 688:20]
  assign _GEN_92 = exception ? _GEN_74 : reg_mstatus_mie; // @[CSR.scala 688:20]
  assign _GEN_95 = io_rw_addr[10] ? ~_T_400 : ~_T_374; // @[CSR.scala 745:53]
  assign _GEN_100 = ~io_rw_addr[9] | _GEN_84; // @[CSR.scala 739:52]
  assign _GEN_101 = io_rw_addr[9] ? _GEN_85 : 2'h0; // @[CSR.scala 739:52]
  assign _GEN_103 = io_rw_addr[9] ? _GEN_95 : ~_T_450; // @[CSR.scala 739:52]
  assign _GEN_110 = insn_ret ? _GEN_101 : _GEN_85; // @[CSR.scala 738:19]
  assign _GEN_112 = insn_ret ? {{24'd0}, _GEN_103} : tvec; // @[CSR.scala 738:19]
  assign _GEN_117 = insn_cease | _T_1579; // @[Reg.scala 28:19]
  assign _T_1581 = _T_552 ? _T_366 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1582 = _T_553 ? _T_370 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1583 = _T_554 ? reg_misa : 64'h0; // @[Mux.scala 27:72]
  assign _T_1584 = _T_555 ? read_mstatus : 64'h0; // @[Mux.scala 27:72]
  assign _T_1585 = _T_556 ? read_mtvec : 64'h0; // @[Mux.scala 27:72]
  assign _T_1586 = _T_557 ? read_mip : 16'h0; // @[Mux.scala 27:72]
  assign _T_1587 = _T_558 ? reg_mie : 64'h0; // @[Mux.scala 27:72]
  assign _T_1588 = _T_559 ? reg_mscratch : 64'h0; // @[Mux.scala 27:72]
  assign _T_1589 = _T_560 ? _T_379 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1590 = _T_561 ? _T_383 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1591 = _T_562 ? reg_mcause : 64'h0; // @[Mux.scala 27:72]
  assign _T_1592 = _T_563 & io_hartid; // @[Mux.scala 27:72]
  assign _T_1593 = _T_564 ? _T_396 : 32'h0; // @[Mux.scala 27:72]
  assign _T_1594 = _T_565 ? _T_405 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1595 = _T_566 ? reg_dscratch : 64'h0; // @[Mux.scala 27:72]
  assign _T_1596 = _T_567 ? reg_fflags : 5'h0; // @[Mux.scala 27:72]
  assign _T_1597 = _T_568 ? reg_frm : 3'h0; // @[Mux.scala 27:72]
  assign _T_1598 = _T_569 ? read_fcsr : 8'h0; // @[Mux.scala 27:72]
  assign _T_1599 = _T_570 ? _T_53 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1600 = _T_571 ? _T_45 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1688 = _T_659 ? read_mcounteren : 32'h0; // @[Mux.scala 27:72]
  assign _T_1689 = _T_660 ? _T_53 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1690 = _T_661 ? _T_45 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1691 = _T_662 ? _T_439[63:0] : 64'h0; // @[Mux.scala 27:72]
  assign _T_1692 = _T_663 ? _T_407 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1693 = _T_664 ? _T_406 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1694 = _T_665 ? reg_sscratch : 64'h0; // @[Mux.scala 27:72]
  assign _T_1695 = _T_666 ? reg_scause : 64'h0; // @[Mux.scala 27:72]
  assign _T_1696 = _T_667 ? _T_444 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1697 = _T_668 ? _T_446 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1698 = _T_669 ? _T_455 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1699 = _T_670 ? read_stvec : 64'h0; // @[Mux.scala 27:72]
  assign _T_1700 = _T_671 ? read_scounteren : 32'h0; // @[Mux.scala 27:72]
  assign _T_1701 = _T_672 ? read_mideleg : 64'h0; // @[Mux.scala 27:72]
  assign _T_1702 = _T_673 ? read_medeleg : 64'h0; // @[Mux.scala 27:72]
  assign _T_1703 = _T_674 ? _T_503 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1705 = _T_676 ? reg_pmp_0_addr : 30'h0; // @[Mux.scala 27:72]
  assign _T_1706 = _T_677 ? reg_pmp_1_addr : 30'h0; // @[Mux.scala 27:72]
  assign _T_1707 = _T_678 ? reg_pmp_2_addr : 30'h0; // @[Mux.scala 27:72]
  assign _T_1708 = _T_679 ? reg_pmp_3_addr : 30'h0; // @[Mux.scala 27:72]
  assign _T_1709 = _T_680 ? reg_pmp_4_addr : 30'h0; // @[Mux.scala 27:72]
  assign _T_1710 = _T_681 ? reg_pmp_5_addr : 30'h0; // @[Mux.scala 27:72]
  assign _T_1711 = _T_682 ? reg_pmp_6_addr : 30'h0; // @[Mux.scala 27:72]
  assign _T_1712 = _T_683 ? reg_pmp_7_addr : 30'h0; // @[Mux.scala 27:72]
  assign _T_1721 = _T_692 ? reg_custom_0 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1722 = _T_693 ? 64'h1 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1724 = _T_695 ? 64'h20181004 : 64'h0; // @[Mux.scala 27:72]
  assign _T_1726 = _T_1581 | _T_1582; // @[Mux.scala 27:72]
  assign _T_1727 = _T_1726 | _T_1583; // @[Mux.scala 27:72]
  assign _T_1728 = _T_1727 | _T_1584; // @[Mux.scala 27:72]
  assign _T_1729 = _T_1728 | _T_1585; // @[Mux.scala 27:72]
  assign _GEN_502 = {{48'd0}, _T_1586}; // @[Mux.scala 27:72]
  assign _T_1730 = _T_1729 | _GEN_502; // @[Mux.scala 27:72]
  assign _T_1731 = _T_1730 | _T_1587; // @[Mux.scala 27:72]
  assign _T_1732 = _T_1731 | _T_1588; // @[Mux.scala 27:72]
  assign _T_1733 = _T_1732 | _T_1589; // @[Mux.scala 27:72]
  assign _T_1734 = _T_1733 | _T_1590; // @[Mux.scala 27:72]
  assign _T_1735 = _T_1734 | _T_1591; // @[Mux.scala 27:72]
  assign _GEN_503 = {{63'd0}, _T_1592}; // @[Mux.scala 27:72]
  assign _T_1736 = _T_1735 | _GEN_503; // @[Mux.scala 27:72]
  assign _GEN_504 = {{32'd0}, _T_1593}; // @[Mux.scala 27:72]
  assign _T_1737 = _T_1736 | _GEN_504; // @[Mux.scala 27:72]
  assign _T_1738 = _T_1737 | _T_1594; // @[Mux.scala 27:72]
  assign _T_1739 = _T_1738 | _T_1595; // @[Mux.scala 27:72]
  assign _GEN_505 = {{59'd0}, _T_1596}; // @[Mux.scala 27:72]
  assign _T_1740 = _T_1739 | _GEN_505; // @[Mux.scala 27:72]
  assign _GEN_506 = {{61'd0}, _T_1597}; // @[Mux.scala 27:72]
  assign _T_1741 = _T_1740 | _GEN_506; // @[Mux.scala 27:72]
  assign _GEN_507 = {{56'd0}, _T_1598}; // @[Mux.scala 27:72]
  assign _T_1742 = _T_1741 | _GEN_507; // @[Mux.scala 27:72]
  assign _T_1743 = _T_1742 | _T_1599; // @[Mux.scala 27:72]
  assign _T_1744 = _T_1743 | _T_1600; // @[Mux.scala 27:72]
  assign _GEN_508 = {{32'd0}, _T_1688}; // @[Mux.scala 27:72]
  assign _T_1832 = _T_1744 | _GEN_508; // @[Mux.scala 27:72]
  assign _T_1833 = _T_1832 | _T_1689; // @[Mux.scala 27:72]
  assign _T_1834 = _T_1833 | _T_1690; // @[Mux.scala 27:72]
  assign _T_1835 = _T_1834 | _T_1691; // @[Mux.scala 27:72]
  assign _T_1836 = _T_1835 | _T_1692; // @[Mux.scala 27:72]
  assign _T_1837 = _T_1836 | _T_1693; // @[Mux.scala 27:72]
  assign _T_1838 = _T_1837 | _T_1694; // @[Mux.scala 27:72]
  assign _T_1839 = _T_1838 | _T_1695; // @[Mux.scala 27:72]
  assign _T_1840 = _T_1839 | _T_1696; // @[Mux.scala 27:72]
  assign _T_1841 = _T_1840 | _T_1697; // @[Mux.scala 27:72]
  assign _T_1842 = _T_1841 | _T_1698; // @[Mux.scala 27:72]
  assign _T_1843 = _T_1842 | _T_1699; // @[Mux.scala 27:72]
  assign _GEN_509 = {{32'd0}, _T_1700}; // @[Mux.scala 27:72]
  assign _T_1844 = _T_1843 | _GEN_509; // @[Mux.scala 27:72]
  assign _T_1845 = _T_1844 | _T_1701; // @[Mux.scala 27:72]
  assign _T_1846 = _T_1845 | _T_1702; // @[Mux.scala 27:72]
  assign _T_1847 = _T_1846 | _T_1703; // @[Mux.scala 27:72]
  assign _GEN_510 = {{34'd0}, _T_1705}; // @[Mux.scala 27:72]
  assign _T_1849 = _T_1847 | _GEN_510; // @[Mux.scala 27:72]
  assign _GEN_511 = {{34'd0}, _T_1706}; // @[Mux.scala 27:72]
  assign _T_1850 = _T_1849 | _GEN_511; // @[Mux.scala 27:72]
  assign _GEN_512 = {{34'd0}, _T_1707}; // @[Mux.scala 27:72]
  assign _T_1851 = _T_1850 | _GEN_512; // @[Mux.scala 27:72]
  assign _GEN_513 = {{34'd0}, _T_1708}; // @[Mux.scala 27:72]
  assign _T_1852 = _T_1851 | _GEN_513; // @[Mux.scala 27:72]
  assign _GEN_514 = {{34'd0}, _T_1709}; // @[Mux.scala 27:72]
  assign _T_1853 = _T_1852 | _GEN_514; // @[Mux.scala 27:72]
  assign _GEN_515 = {{34'd0}, _T_1710}; // @[Mux.scala 27:72]
  assign _T_1854 = _T_1853 | _GEN_515; // @[Mux.scala 27:72]
  assign _GEN_516 = {{34'd0}, _T_1711}; // @[Mux.scala 27:72]
  assign _T_1855 = _T_1854 | _GEN_516; // @[Mux.scala 27:72]
  assign _GEN_517 = {{34'd0}, _T_1712}; // @[Mux.scala 27:72]
  assign _T_1856 = _T_1855 | _GEN_517; // @[Mux.scala 27:72]
  assign _T_1865 = _T_1856 | _T_1721; // @[Mux.scala 27:72]
  assign _T_1866 = _T_1865 | _T_1722; // @[Mux.scala 27:72]
  assign _T_1872 = io_rw_cmd == 3'h5; // @[package.scala 15:47]
  assign _T_1873 = io_rw_cmd == 3'h6; // @[package.scala 15:47]
  assign _T_1874 = io_rw_cmd == 3'h7; // @[package.scala 15:47]
  assign _T_3610 = reg_fflags | io_fcsr_flags_bits; // @[CSR.scala 798:30]
  assign _GEN_118 = io_fcsr_flags_valid ? _T_3610 : reg_fflags; // @[CSR.scala 797:30]
  assign _T_3614 = _T_1873 | _T_1874; // @[package.scala 64:59]
  assign csr_wen = _T_3614 | _T_1872; // @[package.scala 64:59]
  assign _T_3628 = {{39'd0}, wdata};
  assign _T_3660 = _T_3628[12:11] == 2'h2; // @[CSR.scala 1073:35]
  assign _T_3662 = |_T_3628[14:13]; // @[CSR.scala 1094:73]
  assign _GEN_124 = _T_555 ? {{1'd0}, _T_3628[8]} : _GEN_110; // @[CSR.scala 812:39]
  assign _T_3670 = ~io_pc[1] | wdata[2]; // @[CSR.scala 841:43]
  assign _T_3673 = {~wdata[5], 3'h0}; // @[CSR.scala 843:38]
  assign _GEN_518 = {{60'd0}, _T_3673}; // @[CSR.scala 843:32]
  assign _T_3674 = ~wdata | _GEN_518; // @[CSR.scala 843:32]
  assign _T_3676 = ~_T_3674 & 64'h102d; // @[CSR.scala 843:55]
  assign _T_3678 = reg_misa & 64'hffffffffffffefd2; // @[CSR.scala 843:73]
  assign _T_3679 = _T_3676 | _T_3678; // @[CSR.scala 843:62]
  assign _T_3694 = {4'h0,2'h0,reg_mip_seip,1'h0,2'h0,reg_mip_stip,1'h0,2'h0,reg_mip_ssip,1'h0}; // @[CSR.scala 851:59]
  assign _T_3696 = io_rw_cmd[1] ? _T_3694 : 16'h0; // @[CSR.scala 1069:9]
  assign _GEN_519 = {{48'd0}, _T_3696}; // @[CSR.scala 1069:34]
  assign _T_3697 = _GEN_519 | io_rw_wdata; // @[CSR.scala 1069:34]
  assign _T_3702 = _T_3697 & ~_T_701; // @[CSR.scala 1069:43]
  assign _T_3721 = wdata & 64'haaa; // @[CSR.scala 858:59]
  assign _T_3723 = ~wdata | 64'h1; // @[CSR.scala 1090:31]
  assign _GEN_140 = _T_560 ? ~_T_3723 : {{24'd0}, _GEN_87}; // @[CSR.scala 859:40]
  assign _GEN_142 = _T_556 ? wdata : {{32'd0}, reg_mtvec}; // @[CSR.scala 862:40]
  assign _T_3725 = wdata & 64'h800000000000000f; // @[CSR.scala 863:62]
  assign _GEN_145 = _T_570 ? wdata : {{57'd0}, _T_48}; // @[CSR.scala 1087:31]
  assign _GEN_147 = _T_571 ? wdata : {{57'd0}, _T_40}; // @[CSR.scala 1087:31]
  assign _GEN_150 = _T_567 ? wdata : {{59'd0}, _GEN_118}; // @[CSR.scala 876:40]
  assign _GEN_152 = _T_568 ? wdata : {{61'd0}, reg_frm}; // @[CSR.scala 877:40]
  assign _GEN_154 = _T_569 ? wdata : _GEN_150; // @[CSR.scala 878:38]
  assign _GEN_155 = _T_569 ? {{5'd0}, wdata[63:5]} : _GEN_152; // @[CSR.scala 878:38]
  assign _T_3748 = wdata[1:0] == 2'h2; // @[CSR.scala 1073:35]
  assign _GEN_161 = _T_565 ? ~_T_3723 : {{24'd0}, _GEN_76}; // @[CSR.scala 893:42]
  assign _GEN_165 = _T_662 ? {{1'd0}, _T_3628[8]} : _GEN_124; // @[CSR.scala 897:41]
  assign _T_3790 = _GEN_493 & ~read_mideleg; // @[CSR.scala 910:52]
  assign _T_3791 = wdata & read_mideleg; // @[CSR.scala 910:78]
  assign _T_3792 = _T_3790 | _T_3791; // @[CSR.scala 910:69]
  assign _T_3816 = wdata[63:60] == 4'h0; // @[package.scala 15:47]
  assign _T_3817 = wdata[63:60] == 4'h8; // @[package.scala 15:47]
  assign _T_3818 = _T_3816 | _T_3817; // @[package.scala 64:59]
  assign _T_3819 = wdata[63:60] & 4'h8; // @[CSR.scala 918:44]
  assign _T_3822 = reg_mie & ~read_mideleg; // @[CSR.scala 924:64]
  assign _T_3824 = _T_3822 | _T_3791; // @[CSR.scala 924:81]
  assign _GEN_177 = _T_669 ? ~_T_3723 : {{24'd0}, _GEN_80}; // @[CSR.scala 926:42]
  assign _GEN_178 = _T_670 ? wdata : {{25'd0}, reg_stvec}; // @[CSR.scala 927:42]
  assign _T_3828 = wdata & 64'h800000000000001f; // @[CSR.scala 928:64]
  assign _GEN_183 = _T_671 ? wdata : {{32'd0}, reg_scounteren}; // @[CSR.scala 932:44]
  assign _GEN_184 = _T_659 ? wdata : {{32'd0}, reg_mcounteren}; // @[CSR.scala 935:44]
  assign _T_3832 = ~reg_bp_0_control_dmode | reg_debug; // @[CSR.scala 941:55]
  assign _GEN_186 = _T_553 ? wdata : {{25'd0}, reg_bp_0_address}; // @[CSR.scala 942:44]
  assign _T_3866 = io_rw_cmd[1] ? _T_366 : 64'h0; // @[CSR.scala 1069:9]
  assign _T_3867 = _T_3866 | io_rw_wdata; // @[CSR.scala 1069:34]
  assign _T_3872 = _T_3867 & ~_T_701; // @[CSR.scala 1069:43]
  assign _T_3890 = _T_3872[59] & reg_debug; // @[CSR.scala 951:38]
  assign _GEN_187 = _T_3890 & _T_3872[12]; // @[CSR.scala 953:51]
  assign _GEN_203 = _T_3832 ? _GEN_186 : {{25'd0}, reg_bp_0_address}; // @[CSR.scala 941:70]
  assign _T_3975 = _T_674 & ~reg_pmp_0_cfg_l; // @[CSR.scala 961:57]
  assign _T_3985 = wdata[1] & wdata[0]; // @[CSR.scala 965:31]
  assign _T_3989 = ~reg_pmp_1_cfg_a[1] & reg_pmp_1_cfg_a[0]; // @[PMP.scala 49:20]
  assign _T_3990 = reg_pmp_1_cfg_l & _T_3989; // @[PMP.scala 51:62]
  assign _T_3991 = reg_pmp_0_cfg_l | _T_3990; // @[PMP.scala 51:44]
  assign _T_3993 = _T_676 & ~_T_3991; // @[CSR.scala 970:45]
  assign _GEN_258 = _T_3993 ? wdata : {{34'd0}, reg_pmp_0_addr}; // @[CSR.scala 970:71]
  assign _T_3995 = _T_674 & ~reg_pmp_1_cfg_l; // @[CSR.scala 961:57]
  assign _T_4005 = wdata[9] & wdata[8]; // @[CSR.scala 965:31]
  assign _T_4009 = ~reg_pmp_2_cfg_a[1] & reg_pmp_2_cfg_a[0]; // @[PMP.scala 49:20]
  assign _T_4010 = reg_pmp_2_cfg_l & _T_4009; // @[PMP.scala 51:62]
  assign _T_4011 = reg_pmp_1_cfg_l | _T_4010; // @[PMP.scala 51:44]
  assign _T_4013 = _T_677 & ~_T_4011; // @[CSR.scala 970:45]
  assign _GEN_265 = _T_4013 ? wdata : {{34'd0}, reg_pmp_1_addr}; // @[CSR.scala 970:71]
  assign _T_4015 = _T_674 & ~reg_pmp_2_cfg_l; // @[CSR.scala 961:57]
  assign _T_4025 = wdata[17] & wdata[16]; // @[CSR.scala 965:31]
  assign _T_4029 = ~reg_pmp_3_cfg_a[1] & reg_pmp_3_cfg_a[0]; // @[PMP.scala 49:20]
  assign _T_4030 = reg_pmp_3_cfg_l & _T_4029; // @[PMP.scala 51:62]
  assign _T_4031 = reg_pmp_2_cfg_l | _T_4030; // @[PMP.scala 51:44]
  assign _T_4033 = _T_678 & ~_T_4031; // @[CSR.scala 970:45]
  assign _GEN_272 = _T_4033 ? wdata : {{34'd0}, reg_pmp_2_addr}; // @[CSR.scala 970:71]
  assign _T_4035 = _T_674 & ~reg_pmp_3_cfg_l; // @[CSR.scala 961:57]
  assign _T_4045 = wdata[25] & wdata[24]; // @[CSR.scala 965:31]
  assign _T_4049 = ~reg_pmp_4_cfg_a[1] & reg_pmp_4_cfg_a[0]; // @[PMP.scala 49:20]
  assign _T_4050 = reg_pmp_4_cfg_l & _T_4049; // @[PMP.scala 51:62]
  assign _T_4051 = reg_pmp_3_cfg_l | _T_4050; // @[PMP.scala 51:44]
  assign _T_4053 = _T_679 & ~_T_4051; // @[CSR.scala 970:45]
  assign _GEN_279 = _T_4053 ? wdata : {{34'd0}, reg_pmp_3_addr}; // @[CSR.scala 970:71]
  assign _T_4055 = _T_674 & ~reg_pmp_4_cfg_l; // @[CSR.scala 961:57]
  assign _T_4065 = wdata[33] & wdata[32]; // @[CSR.scala 965:31]
  assign _T_4069 = ~reg_pmp_5_cfg_a[1] & reg_pmp_5_cfg_a[0]; // @[PMP.scala 49:20]
  assign _T_4070 = reg_pmp_5_cfg_l & _T_4069; // @[PMP.scala 51:62]
  assign _T_4071 = reg_pmp_4_cfg_l | _T_4070; // @[PMP.scala 51:44]
  assign _T_4073 = _T_680 & ~_T_4071; // @[CSR.scala 970:45]
  assign _GEN_286 = _T_4073 ? wdata : {{34'd0}, reg_pmp_4_addr}; // @[CSR.scala 970:71]
  assign _T_4075 = _T_674 & ~reg_pmp_5_cfg_l; // @[CSR.scala 961:57]
  assign _T_4085 = wdata[41] & wdata[40]; // @[CSR.scala 965:31]
  assign _T_4089 = ~reg_pmp_6_cfg_a[1] & reg_pmp_6_cfg_a[0]; // @[PMP.scala 49:20]
  assign _T_4090 = reg_pmp_6_cfg_l & _T_4089; // @[PMP.scala 51:62]
  assign _T_4091 = reg_pmp_5_cfg_l | _T_4090; // @[PMP.scala 51:44]
  assign _T_4093 = _T_681 & ~_T_4091; // @[CSR.scala 970:45]
  assign _GEN_293 = _T_4093 ? wdata : {{34'd0}, reg_pmp_5_addr}; // @[CSR.scala 970:71]
  assign _T_4095 = _T_674 & ~reg_pmp_6_cfg_l; // @[CSR.scala 961:57]
  assign _T_4105 = wdata[49] & wdata[48]; // @[CSR.scala 965:31]
  assign _T_4109 = ~reg_pmp_7_cfg_a[1] & reg_pmp_7_cfg_a[0]; // @[PMP.scala 49:20]
  assign _T_4110 = reg_pmp_7_cfg_l & _T_4109; // @[PMP.scala 51:62]
  assign _T_4111 = reg_pmp_6_cfg_l | _T_4110; // @[PMP.scala 51:44]
  assign _T_4113 = _T_682 & ~_T_4111; // @[CSR.scala 970:45]
  assign _GEN_300 = _T_4113 ? wdata : {{34'd0}, reg_pmp_6_addr}; // @[CSR.scala 970:71]
  assign _T_4115 = _T_674 & ~reg_pmp_7_cfg_l; // @[CSR.scala 961:57]
  assign _T_4125 = wdata[57] & wdata[56]; // @[CSR.scala 965:31]
  assign _T_4131 = reg_pmp_7_cfg_l | _T_4110; // @[PMP.scala 51:44]
  assign _T_4133 = _T_683 & ~_T_4131; // @[CSR.scala 970:45]
  assign _GEN_307 = _T_4133 ? wdata : {{34'd0}, reg_pmp_7_addr}; // @[CSR.scala 970:71]
  assign _T_4134 = wdata & 64'h208; // @[CSR.scala 977:23]
  assign _T_4136 = reg_custom_0 & 64'hfffffffffffffdf7; // @[CSR.scala 977:38]
  assign _T_4137 = _T_4134 | _T_4136; // @[CSR.scala 977:31]
  assign _GEN_320 = csr_wen ? _GEN_165 : _GEN_110; // @[CSR.scala 811:18]
  assign _GEN_335 = csr_wen ? _GEN_140 : {{24'd0}, _GEN_87}; // @[CSR.scala 811:18]
  assign _GEN_337 = csr_wen ? _GEN_142 : {{32'd0}, reg_mtvec}; // @[CSR.scala 811:18]
  assign _GEN_340 = csr_wen ? _GEN_145 : {{57'd0}, _T_48}; // @[CSR.scala 811:18]
  assign _GEN_342 = csr_wen ? _GEN_147 : {{57'd0}, _T_40}; // @[CSR.scala 811:18]
  assign _GEN_345 = csr_wen ? _GEN_154 : {{59'd0}, _GEN_118}; // @[CSR.scala 811:18]
  assign _GEN_346 = csr_wen ? _GEN_155 : {{61'd0}, reg_frm}; // @[CSR.scala 811:18]
  assign _GEN_352 = csr_wen ? _GEN_161 : {{24'd0}, _GEN_76}; // @[CSR.scala 811:18]
  assign _GEN_357 = csr_wen ? _GEN_177 : {{24'd0}, _GEN_80}; // @[CSR.scala 811:18]
  assign _GEN_358 = csr_wen ? _GEN_178 : {{25'd0}, reg_stvec}; // @[CSR.scala 811:18]
  assign _GEN_363 = csr_wen ? _GEN_183 : {{32'd0}, reg_scounteren}; // @[CSR.scala 811:18]
  assign _GEN_364 = csr_wen ? _GEN_184 : {{32'd0}, reg_mcounteren}; // @[CSR.scala 811:18]
  assign _GEN_366 = csr_wen ? _GEN_203 : {{25'd0}, reg_bp_0_address}; // @[CSR.scala 811:18]
  assign _GEN_404 = csr_wen ? _GEN_258 : {{34'd0}, reg_pmp_0_addr}; // @[CSR.scala 811:18]
  assign _GEN_411 = csr_wen ? _GEN_265 : {{34'd0}, reg_pmp_1_addr}; // @[CSR.scala 811:18]
  assign _GEN_418 = csr_wen ? _GEN_272 : {{34'd0}, reg_pmp_2_addr}; // @[CSR.scala 811:18]
  assign _GEN_425 = csr_wen ? _GEN_279 : {{34'd0}, reg_pmp_3_addr}; // @[CSR.scala 811:18]
  assign _GEN_432 = csr_wen ? _GEN_286 : {{34'd0}, reg_pmp_4_addr}; // @[CSR.scala 811:18]
  assign _GEN_439 = csr_wen ? _GEN_293 : {{34'd0}, reg_pmp_5_addr}; // @[CSR.scala 811:18]
  assign _GEN_446 = csr_wen ? _GEN_300 : {{34'd0}, reg_pmp_6_addr}; // @[CSR.scala 811:18]
  assign _GEN_453 = csr_wen ? _GEN_307 : {{34'd0}, reg_pmp_7_addr}; // @[CSR.scala 811:18]
  assign _T_4163 = io_retire > 1'h0; // @[CSR.scala 1048:26]
  assign io_rw_rdata = _T_1866 | _T_1724; // @[CSR.scala 769:15]
  assign io_decode_0_fp_illegal = _T_782 | ~reg_misa[5]; // @[CSR.scala 616:23]
  assign io_decode_0_fp_csr = _T_790 == 12'h0; // @[CSR.scala 618:19]
  assign io_decode_0_read_illegal = _T_1111 | _T_1114; // @[CSR.scala 620:25]
  assign io_decode_0_write_illegal = &io_decode_0_csr[11:10]; // @[CSR.scala 627:26]
  assign io_decode_0_write_flush = ~_T_1124; // @[CSR.scala 628:24]
  assign io_decode_0_system_illegal = _T_1138 | _T_1140; // @[CSR.scala 629:27]
  assign io_csr_stall = reg_wfi | io_status_cease; // @[CSR.scala 759:16]
  assign io_eret = _T_1197 | insn_ret; // @[CSR.scala 661:11]
  assign io_singleStep = reg_dcsr_step & ~reg_debug; // @[CSR.scala 662:17]
  assign io_status_debug = reg_debug; // @[CSR.scala 663:13 CSR.scala 665:19]
  assign io_status_cease = _T_1579; // @[CSR.scala 663:13 CSR.scala 760:19]
  assign io_status_wfi = reg_wfi; // @[CSR.scala 663:13 CSR.scala 761:17]
  assign io_status_isa = reg_misa[31:0]; // @[CSR.scala 663:13 CSR.scala 666:17]
  assign io_status_dprv = _T_1196; // @[CSR.scala 663:13 CSR.scala 669:18]
  assign io_status_prv = reg_mstatus_prv; // @[CSR.scala 663:13]
  assign io_status_sd = _T_1190 | _T_1191; // @[CSR.scala 663:13 CSR.scala 664:16]
  assign io_status_zero2 = 27'h0; // @[CSR.scala 663:13]
  assign io_status_sxl = 2'h2; // @[CSR.scala 663:13 CSR.scala 668:17]
  assign io_status_uxl = 2'h2; // @[CSR.scala 663:13 CSR.scala 667:17]
  assign io_status_sd_rv32 = 1'h0; // @[CSR.scala 663:13]
  assign io_status_zero1 = 8'h0; // @[CSR.scala 663:13]
  assign io_status_tsr = reg_mstatus_tsr; // @[CSR.scala 663:13]
  assign io_status_tw = reg_mstatus_tw; // @[CSR.scala 663:13]
  assign io_status_tvm = reg_mstatus_tvm; // @[CSR.scala 663:13]
  assign io_status_mxr = reg_mstatus_mxr; // @[CSR.scala 663:13]
  assign io_status_sum = reg_mstatus_sum; // @[CSR.scala 663:13]
  assign io_status_mprv = reg_mstatus_mprv; // @[CSR.scala 663:13]
  assign io_status_xs = 2'h0; // @[CSR.scala 663:13]
  assign io_status_fs = reg_mstatus_fs; // @[CSR.scala 663:13]
  assign io_status_mpp = reg_mstatus_mpp; // @[CSR.scala 663:13]
  assign io_status_vs = 2'h0; // @[CSR.scala 663:13]
  assign io_status_spp = reg_mstatus_spp; // @[CSR.scala 663:13]
  assign io_status_mpie = reg_mstatus_mpie; // @[CSR.scala 663:13]
  assign io_status_hpie = 1'h0; // @[CSR.scala 663:13]
  assign io_status_spie = reg_mstatus_spie; // @[CSR.scala 663:13]
  assign io_status_upie = 1'h0; // @[CSR.scala 663:13]
  assign io_status_mie = reg_mstatus_mie; // @[CSR.scala 663:13]
  assign io_status_hie = 1'h0; // @[CSR.scala 663:13]
  assign io_status_sie = reg_mstatus_sie; // @[CSR.scala 663:13]
  assign io_status_uie = 1'h0; // @[CSR.scala 663:13]
  assign io_ptbr_mode = reg_satp_mode; // @[CSR.scala 660:11]
  assign io_ptbr_ppn = reg_satp_ppn; // @[CSR.scala 660:11]
  assign io_evec = _GEN_112[39:0]; // @[CSR.scala 659:11 CSR.scala 744:15 CSR.scala 748:15 CSR.scala 754:15]
  assign io_time = {_T_49,_T_47}; // @[CSR.scala 758:11]
  assign io_fcsr_rm = reg_frm; // @[CSR.scala 796:14]
  assign io_interrupt = _T_232 & ~_T_233; // @[CSR.scala 439:16]
  assign io_interrupt_cause = 64'h8000000000000000 + _GEN_494; // @[CSR.scala 440:22]
  assign io_bp_0_control_action = reg_bp_0_control_action; // @[CSR.scala 441:9]
  assign io_bp_0_control_tmatch = reg_bp_0_control_tmatch; // @[CSR.scala 441:9]
  assign io_bp_0_control_m = reg_bp_0_control_m; // @[CSR.scala 441:9]
  assign io_bp_0_control_s = reg_bp_0_control_s; // @[CSR.scala 441:9]
  assign io_bp_0_control_u = reg_bp_0_control_u; // @[CSR.scala 441:9]
  assign io_bp_0_control_x = reg_bp_0_control_x; // @[CSR.scala 441:9]
  assign io_bp_0_control_w = reg_bp_0_control_w; // @[CSR.scala 441:9]
  assign io_bp_0_control_r = reg_bp_0_control_r; // @[CSR.scala 441:9]
  assign io_bp_0_address = reg_bp_0_address; // @[CSR.scala 441:9]
  assign io_pmp_0_cfg_l = reg_pmp_0_cfg_l; // @[CSR.scala 442:10]
  assign io_pmp_0_cfg_a = reg_pmp_0_cfg_a; // @[CSR.scala 442:10]
  assign io_pmp_0_cfg_x = reg_pmp_0_cfg_x; // @[CSR.scala 442:10]
  assign io_pmp_0_cfg_w = reg_pmp_0_cfg_w; // @[CSR.scala 442:10]
  assign io_pmp_0_cfg_r = reg_pmp_0_cfg_r; // @[CSR.scala 442:10]
  assign io_pmp_0_addr = reg_pmp_0_addr; // @[CSR.scala 442:10]
  assign io_pmp_0_mask = _T_244[31:0]; // @[CSR.scala 442:10]
  assign io_pmp_1_cfg_l = reg_pmp_1_cfg_l; // @[CSR.scala 442:10]
  assign io_pmp_1_cfg_a = reg_pmp_1_cfg_a; // @[CSR.scala 442:10]
  assign io_pmp_1_cfg_x = reg_pmp_1_cfg_x; // @[CSR.scala 442:10]
  assign io_pmp_1_cfg_w = reg_pmp_1_cfg_w; // @[CSR.scala 442:10]
  assign io_pmp_1_cfg_r = reg_pmp_1_cfg_r; // @[CSR.scala 442:10]
  assign io_pmp_1_addr = reg_pmp_1_addr; // @[CSR.scala 442:10]
  assign io_pmp_1_mask = _T_253[31:0]; // @[CSR.scala 442:10]
  assign io_pmp_2_cfg_l = reg_pmp_2_cfg_l; // @[CSR.scala 442:10]
  assign io_pmp_2_cfg_a = reg_pmp_2_cfg_a; // @[CSR.scala 442:10]
  assign io_pmp_2_cfg_x = reg_pmp_2_cfg_x; // @[CSR.scala 442:10]
  assign io_pmp_2_cfg_w = reg_pmp_2_cfg_w; // @[CSR.scala 442:10]
  assign io_pmp_2_cfg_r = reg_pmp_2_cfg_r; // @[CSR.scala 442:10]
  assign io_pmp_2_addr = reg_pmp_2_addr; // @[CSR.scala 442:10]
  assign io_pmp_2_mask = _T_262[31:0]; // @[CSR.scala 442:10]
  assign io_pmp_3_cfg_l = reg_pmp_3_cfg_l; // @[CSR.scala 442:10]
  assign io_pmp_3_cfg_a = reg_pmp_3_cfg_a; // @[CSR.scala 442:10]
  assign io_pmp_3_cfg_x = reg_pmp_3_cfg_x; // @[CSR.scala 442:10]
  assign io_pmp_3_cfg_w = reg_pmp_3_cfg_w; // @[CSR.scala 442:10]
  assign io_pmp_3_cfg_r = reg_pmp_3_cfg_r; // @[CSR.scala 442:10]
  assign io_pmp_3_addr = reg_pmp_3_addr; // @[CSR.scala 442:10]
  assign io_pmp_3_mask = _T_271[31:0]; // @[CSR.scala 442:10]
  assign io_pmp_4_cfg_l = reg_pmp_4_cfg_l; // @[CSR.scala 442:10]
  assign io_pmp_4_cfg_a = reg_pmp_4_cfg_a; // @[CSR.scala 442:10]
  assign io_pmp_4_cfg_x = reg_pmp_4_cfg_x; // @[CSR.scala 442:10]
  assign io_pmp_4_cfg_w = reg_pmp_4_cfg_w; // @[CSR.scala 442:10]
  assign io_pmp_4_cfg_r = reg_pmp_4_cfg_r; // @[CSR.scala 442:10]
  assign io_pmp_4_addr = reg_pmp_4_addr; // @[CSR.scala 442:10]
  assign io_pmp_4_mask = _T_280[31:0]; // @[CSR.scala 442:10]
  assign io_pmp_5_cfg_l = reg_pmp_5_cfg_l; // @[CSR.scala 442:10]
  assign io_pmp_5_cfg_a = reg_pmp_5_cfg_a; // @[CSR.scala 442:10]
  assign io_pmp_5_cfg_x = reg_pmp_5_cfg_x; // @[CSR.scala 442:10]
  assign io_pmp_5_cfg_w = reg_pmp_5_cfg_w; // @[CSR.scala 442:10]
  assign io_pmp_5_cfg_r = reg_pmp_5_cfg_r; // @[CSR.scala 442:10]
  assign io_pmp_5_addr = reg_pmp_5_addr; // @[CSR.scala 442:10]
  assign io_pmp_5_mask = _T_289[31:0]; // @[CSR.scala 442:10]
  assign io_pmp_6_cfg_l = reg_pmp_6_cfg_l; // @[CSR.scala 442:10]
  assign io_pmp_6_cfg_a = reg_pmp_6_cfg_a; // @[CSR.scala 442:10]
  assign io_pmp_6_cfg_x = reg_pmp_6_cfg_x; // @[CSR.scala 442:10]
  assign io_pmp_6_cfg_w = reg_pmp_6_cfg_w; // @[CSR.scala 442:10]
  assign io_pmp_6_cfg_r = reg_pmp_6_cfg_r; // @[CSR.scala 442:10]
  assign io_pmp_6_addr = reg_pmp_6_addr; // @[CSR.scala 442:10]
  assign io_pmp_6_mask = _T_298[31:0]; // @[CSR.scala 442:10]
  assign io_pmp_7_cfg_l = reg_pmp_7_cfg_l; // @[CSR.scala 442:10]
  assign io_pmp_7_cfg_a = reg_pmp_7_cfg_a; // @[CSR.scala 442:10]
  assign io_pmp_7_cfg_x = reg_pmp_7_cfg_x; // @[CSR.scala 442:10]
  assign io_pmp_7_cfg_w = reg_pmp_7_cfg_w; // @[CSR.scala 442:10]
  assign io_pmp_7_cfg_r = reg_pmp_7_cfg_r; // @[CSR.scala 442:10]
  assign io_pmp_7_addr = reg_pmp_7_addr; // @[CSR.scala 442:10]
  assign io_pmp_7_mask = _T_307[31:0]; // @[CSR.scala 442:10]
  assign io_trace_0_valid = _T_4163 | io_trace_0_exception; // @[CSR.scala 1048:13]
  assign io_trace_0_iaddr = io_pc; // @[CSR.scala 1050:13]
  assign io_trace_0_insn = io_inst_0; // @[CSR.scala 1049:12]
  assign io_trace_0_exception = _T_1197 | io_exception; // @[CSR.scala 1047:17]
  assign io_customCSRs_0_value = reg_custom_0; // @[CSR.scala 766:14]
  assign CSRFile_cov_read_addr = CSRFile_state;
  assign CSRFile_cov_read_data = CSRFile_cov[CSRFile_cov_read_addr]; // @[Coverage map for CSRFile]
  assign CSRFile_cov_write_data = 1'h1;
  assign CSRFile_cov_write_addr = CSRFile_state;
  assign CSRFile_cov_write_mask = 1'h1;
  assign CSRFile_cov_write_en = 1'h1;
  assign reg_dcsr_ebreaku_shl = {reg_dcsr_ebreaku, 1'h0};
  assign reg_dcsr_ebreaku_pad = {18'h0,reg_dcsr_ebreaku_shl};
  assign reg_pmp_3_cfg_l_shl = {reg_pmp_3_cfg_l, 2'h0};
  assign reg_pmp_3_cfg_l_pad = {17'h0,reg_pmp_3_cfg_l_shl};
  assign reg_pmp_5_cfg_l_shl = {reg_pmp_5_cfg_l, 7'h0};
  assign reg_pmp_5_cfg_l_pad = {12'h0,reg_pmp_5_cfg_l_shl};
  assign reg_dcsr_ebreaks_shl = {reg_dcsr_ebreaks, 13'h0};
  assign reg_dcsr_ebreaks_pad = {6'h0,reg_dcsr_ebreaks_shl};
  assign reg_pmp_6_cfg_l_shl = {reg_pmp_6_cfg_l, 14'h0};
  assign reg_pmp_6_cfg_l_pad = {5'h0,reg_pmp_6_cfg_l_shl};
  assign reg_mip_ssip_shl = {reg_mip_ssip, 10'h0};
  assign reg_mip_ssip_pad = {9'h0,reg_mip_ssip_shl};
  assign reg_mip_seip_shl = {reg_mip_seip, 6'h0};
  assign reg_mip_seip_pad = {13'h0,reg_mip_seip_shl};
  assign reg_pmp_7_cfg_l_shl = {reg_pmp_7_cfg_l, 7'h0};
  assign reg_pmp_7_cfg_l_pad = {12'h0,reg_pmp_7_cfg_l_shl};
  assign reg_dcsr_ebreakm_shl = {reg_dcsr_ebreakm, 19'h0};
  assign reg_dcsr_ebreakm_pad = reg_dcsr_ebreakm_shl;
  assign reg_mstatus_spp_shl = {reg_mstatus_spp, 4'h0};
  assign reg_mstatus_spp_pad = {15'h0,reg_mstatus_spp_shl};
  assign reg_debug_shl = {reg_debug, 14'h0};
  assign reg_debug_pad = {5'h0,reg_debug_shl};
  assign reg_pmp_0_cfg_l_shl = {reg_pmp_0_cfg_l, 19'h0};
  assign reg_pmp_0_cfg_l_pad = reg_pmp_0_cfg_l_shl;
  assign reg_mstatus_mprv_shl = {reg_mstatus_mprv, 12'h0};
  assign reg_mstatus_mprv_pad = {7'h0,reg_mstatus_mprv_shl};
  assign reg_pmp_4_cfg_l_shl = {reg_pmp_4_cfg_l, 19'h0};
  assign reg_pmp_4_cfg_l_pad = reg_pmp_4_cfg_l_shl;
  assign reg_singleStepped_shl = {reg_singleStepped, 19'h0};
  assign reg_singleStepped_pad = reg_singleStepped_shl;
  assign reg_mstatus_mie_shl = {reg_mstatus_mie, 4'h0};
  assign reg_mstatus_mie_pad = {15'h0,reg_mstatus_mie_shl};
  assign reg_pmp_1_cfg_l_shl = {reg_pmp_1_cfg_l, 19'h0};
  assign reg_pmp_1_cfg_l_pad = reg_pmp_1_cfg_l_shl;
  assign reg_pmp_7_cfg_a_shl = {reg_pmp_7_cfg_a, 7'h0};
  assign reg_pmp_7_cfg_a_pad = {11'h0,reg_pmp_7_cfg_a_shl};
  assign reg_bp_0_control_dmode_shl = {reg_bp_0_control_dmode, 1'h0};
  assign reg_bp_0_control_dmode_pad = {18'h0,reg_bp_0_control_dmode_shl};
  assign reg_mip_stip_shl = {reg_mip_stip, 11'h0};
  assign reg_mip_stip_pad = {8'h0,reg_mip_stip_shl};
  assign reg_mstatus_sie_shl = {reg_mstatus_sie, 15'h0};
  assign reg_mstatus_sie_pad = {4'h0,reg_mstatus_sie_shl};
  assign reg_pmp_2_cfg_l_shl = {reg_pmp_2_cfg_l, 5'h0};
  assign reg_pmp_2_cfg_l_pad = {14'h0,reg_pmp_2_cfg_l_shl};
  assign reg_mstatus_prv_shl = {reg_mstatus_prv, 2'h0};
  assign reg_mstatus_prv_pad = {16'h0,reg_mstatus_prv_shl};
  assign CSRFile_xor7 = reg_dcsr_ebreaku_pad ^ reg_pmp_3_cfg_l_pad;
  assign CSRFile_xor18 = reg_dcsr_ebreaks_pad ^ reg_pmp_6_cfg_l_pad;
  assign CSRFile_xor8 = reg_pmp_5_cfg_l_pad ^ CSRFile_xor18;
  assign CSRFile_xor3 = CSRFile_xor7 ^ CSRFile_xor8;
  assign CSRFile_xor20 = reg_mip_seip_pad ^ reg_pmp_7_cfg_l_pad;
  assign CSRFile_xor9 = reg_mip_ssip_pad ^ CSRFile_xor20;
  assign CSRFile_xor22 = reg_mstatus_spp_pad ^ reg_debug_pad;
  assign CSRFile_xor10 = reg_dcsr_ebreakm_pad ^ CSRFile_xor22;
  assign CSRFile_xor4 = CSRFile_xor9 ^ CSRFile_xor10;
  assign CSRFile_xor1 = CSRFile_xor3 ^ CSRFile_xor4;
  assign CSRFile_xor24 = reg_mstatus_mprv_pad ^ reg_pmp_4_cfg_l_pad;
  assign CSRFile_xor11 = reg_pmp_0_cfg_l_pad ^ CSRFile_xor24;
  assign CSRFile_xor26 = reg_mstatus_mie_pad ^ reg_pmp_1_cfg_l_pad;
  assign CSRFile_xor12 = reg_singleStepped_pad ^ CSRFile_xor26;
  assign CSRFile_xor5 = CSRFile_xor11 ^ CSRFile_xor12;
  assign CSRFile_xor28 = reg_bp_0_control_dmode_pad ^ reg_mip_stip_pad;
  assign CSRFile_xor13 = reg_pmp_7_cfg_a_pad ^ CSRFile_xor28;
  assign CSRFile_xor30 = reg_pmp_2_cfg_l_pad ^ reg_mstatus_prv_pad;
  assign CSRFile_xor14 = reg_mstatus_sie_pad ^ CSRFile_xor30;
  assign CSRFile_xor6 = CSRFile_xor13 ^ CSRFile_xor14;
  assign CSRFile_xor2 = CSRFile_xor5 ^ CSRFile_xor6;
  assign CSRFile_xor0 = CSRFile_xor1 ^ CSRFile_xor2;
  assign io_covSum = CSRFile_covSum;
  assign stopEn0 = ~_T_1206;
  assign stopEn1 = ~_T_1228;
  assign CSRFile_or0 = stopEn0 | stopEn1;
  assign metaAssert = CSRFile_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_prv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_tsr = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus_tw = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_mstatus_tvm = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_mstatus_mxr = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_mstatus_sum = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_mstatus_mprv = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_mstatus_fs = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_mstatus_mpp = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_mstatus_spp = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_mstatus_spie = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  reg_mstatus_sie = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  reg_dcsr_prv = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  reg_singleStepped = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  reg_dcsr_ebreakm = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  reg_dcsr_ebreaks = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  reg_dcsr_ebreaku = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  reg_debug = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  reg_mideleg = _RAND_20[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  reg_medeleg = _RAND_21[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  reg_dcsr_cause = _RAND_22[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  reg_dcsr_step = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{`RANDOM}};
  reg_dpc = _RAND_24[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{`RANDOM}};
  reg_dscratch = _RAND_25[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  reg_bp_0_control_dmode = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  reg_bp_0_control_action = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  reg_bp_0_control_tmatch = _RAND_28[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  reg_bp_0_control_m = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  reg_bp_0_control_s = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  reg_bp_0_control_u = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  reg_bp_0_control_x = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  reg_bp_0_control_w = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  reg_bp_0_control_r = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{`RANDOM}};
  reg_bp_0_address = _RAND_35[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  reg_pmp_0_cfg_l = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  reg_pmp_0_cfg_a = _RAND_37[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  reg_pmp_0_cfg_x = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  reg_pmp_0_cfg_w = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  reg_pmp_0_cfg_r = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  reg_pmp_0_addr = _RAND_41[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  reg_pmp_1_cfg_l = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  reg_pmp_1_cfg_a = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  reg_pmp_1_cfg_x = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  reg_pmp_1_cfg_w = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  reg_pmp_1_cfg_r = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  reg_pmp_1_addr = _RAND_47[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  reg_pmp_2_cfg_l = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  reg_pmp_2_cfg_a = _RAND_49[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  reg_pmp_2_cfg_x = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  reg_pmp_2_cfg_w = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  reg_pmp_2_cfg_r = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  reg_pmp_2_addr = _RAND_53[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  reg_pmp_3_cfg_l = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  reg_pmp_3_cfg_a = _RAND_55[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  reg_pmp_3_cfg_x = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  reg_pmp_3_cfg_w = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  reg_pmp_3_cfg_r = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  reg_pmp_3_addr = _RAND_59[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  reg_pmp_4_cfg_l = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  reg_pmp_4_cfg_a = _RAND_61[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  reg_pmp_4_cfg_x = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  reg_pmp_4_cfg_w = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  reg_pmp_4_cfg_r = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  reg_pmp_4_addr = _RAND_65[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  reg_pmp_5_cfg_l = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  reg_pmp_5_cfg_a = _RAND_67[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  reg_pmp_5_cfg_x = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  reg_pmp_5_cfg_w = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  reg_pmp_5_cfg_r = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  reg_pmp_5_addr = _RAND_71[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  reg_pmp_6_cfg_l = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  reg_pmp_6_cfg_a = _RAND_73[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  reg_pmp_6_cfg_x = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  reg_pmp_6_cfg_w = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  reg_pmp_6_cfg_r = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  reg_pmp_6_addr = _RAND_77[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  reg_pmp_7_cfg_l = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  reg_pmp_7_cfg_a = _RAND_79[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  reg_pmp_7_cfg_x = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  reg_pmp_7_cfg_w = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  reg_pmp_7_cfg_r = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  reg_pmp_7_addr = _RAND_83[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {2{`RANDOM}};
  reg_mie = _RAND_84[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  reg_mip_seip = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  reg_mip_stip = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  reg_mip_ssip = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {2{`RANDOM}};
  reg_mepc = _RAND_88[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {2{`RANDOM}};
  reg_mcause = _RAND_89[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  reg_mtval = _RAND_90[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {2{`RANDOM}};
  reg_mscratch = _RAND_91[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  reg_mtvec = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  reg_mcounteren = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  reg_scounteren = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {2{`RANDOM}};
  reg_sepc = _RAND_95[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {2{`RANDOM}};
  reg_scause = _RAND_96[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {2{`RANDOM}};
  reg_stval = _RAND_97[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {2{`RANDOM}};
  reg_sscratch = _RAND_98[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {2{`RANDOM}};
  reg_stvec = _RAND_99[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  reg_satp_mode = _RAND_100[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {2{`RANDOM}};
  reg_satp_ppn = _RAND_101[43:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  reg_wfi = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  reg_fflags = _RAND_103[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  reg_frm = _RAND_104[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_39 = _RAND_105[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {2{`RANDOM}};
  _T_41 = _RAND_106[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_47 = _RAND_107[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {2{`RANDOM}};
  _T_49 = _RAND_108[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {2{`RANDOM}};
  reg_misa = _RAND_109[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {2{`RANDOM}};
  reg_custom_0 = _RAND_110[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_1196 = _RAND_111[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_1579 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  CSRFile_state = _RAND_113[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    CSRFile_cov[initvar] = _RAND_114[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  CSRFile_covSum = _RAND_115[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  CSRFile_metaAssert = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      reg_mstatus_prv <= 2'h0;
    end else if (reset) begin
      reg_mstatus_prv <= 2'h3;
    end else if (_T_1) begin
      reg_mstatus_prv <= 2'h0;
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        reg_mstatus_prv <= {{1'd0}, reg_mstatus_spp};
      end else if (io_rw_addr[10]) begin
        reg_mstatus_prv <= reg_dcsr_prv;
      end else begin
        reg_mstatus_prv <= reg_mstatus_mpp;
      end
    end else if (exception) begin
      if (trapToDebug) begin
        if (~reg_debug) begin
          reg_mstatus_prv <= 2'h3;
        end
      end else if (delegate) begin
        reg_mstatus_prv <= 2'h1;
      end else begin
        reg_mstatus_prv <= 2'h3;
      end
    end
    if (metaReset) begin
      reg_mstatus_tsr <= 1'h0;
    end else if (reset) begin
      reg_mstatus_tsr <= 1'h0;
    end else if (csr_wen) begin
      if (_T_555) begin
        reg_mstatus_tsr <= _T_3628[22];
      end
    end
    if (metaReset) begin
      reg_mstatus_tw <= 1'h0;
    end else if (reset) begin
      reg_mstatus_tw <= 1'h0;
    end else if (csr_wen) begin
      if (_T_555) begin
        reg_mstatus_tw <= _T_3628[21];
      end
    end
    if (metaReset) begin
      reg_mstatus_tvm <= 1'h0;
    end else if (reset) begin
      reg_mstatus_tvm <= 1'h0;
    end else if (csr_wen) begin
      if (_T_555) begin
        reg_mstatus_tvm <= _T_3628[20];
      end
    end
    if (metaReset) begin
      reg_mstatus_mxr <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mxr <= 1'h0;
    end else if (csr_wen) begin
      if (_T_662) begin
        reg_mstatus_mxr <= _T_3628[19];
      end else if (_T_555) begin
        reg_mstatus_mxr <= _T_3628[19];
      end
    end
    if (metaReset) begin
      reg_mstatus_sum <= 1'h0;
    end else if (reset) begin
      reg_mstatus_sum <= 1'h0;
    end else if (csr_wen) begin
      if (_T_662) begin
        reg_mstatus_sum <= _T_3628[18];
      end else if (_T_555) begin
        reg_mstatus_sum <= _T_3628[18];
      end
    end
    if (metaReset) begin
      reg_mstatus_mprv <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mprv <= 1'h0;
    end else if (csr_wen) begin
      if (_T_555) begin
        reg_mstatus_mprv <= _T_3628[17];
      end
    end
    if (metaReset) begin
      reg_mstatus_fs <= 2'h0;
    end else if (reset) begin
      reg_mstatus_fs <= 2'h0;
    end else if (csr_wen) begin
      if (_T_662) begin
        if (_T_3662) begin
          reg_mstatus_fs <= 2'h3;
        end else begin
          reg_mstatus_fs <= 2'h0;
        end
      end else if (_T_555) begin
        if (_T_3662) begin
          reg_mstatus_fs <= 2'h3;
        end else begin
          reg_mstatus_fs <= 2'h0;
        end
      end
    end
    if (metaReset) begin
      reg_mstatus_mpp <= 2'h0;
    end else if (reset) begin
      reg_mstatus_mpp <= 2'h3;
    end else if (csr_wen) begin
      if (_T_555) begin
        if (_T_3660) begin
          reg_mstatus_mpp <= 2'h0;
        end else begin
          reg_mstatus_mpp <= _T_3628[12:11];
        end
      end else if (insn_ret) begin
        if (~io_rw_addr[9]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (!(delegate)) begin
                reg_mstatus_mpp <= reg_mstatus_prv;
              end
            end
          end
        end else if (io_rw_addr[10]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (!(delegate)) begin
                reg_mstatus_mpp <= reg_mstatus_prv;
              end
            end
          end
        end else begin
          reg_mstatus_mpp <= 2'h0;
        end
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (!(delegate)) begin
            reg_mstatus_mpp <= reg_mstatus_prv;
          end
        end
      end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        if (exception) begin
          if (!(trapToDebug)) begin
            if (!(delegate)) begin
              reg_mstatus_mpp <= reg_mstatus_prv;
            end
          end
        end
      end else if (io_rw_addr[10]) begin
        reg_mstatus_mpp <= _GEN_91;
      end else begin
        reg_mstatus_mpp <= 2'h0;
      end
    end else begin
      reg_mstatus_mpp <= _GEN_91;
    end
    if (metaReset) begin
      reg_mstatus_spp <= 1'h0;
    end else if (reset) begin
      reg_mstatus_spp <= 1'h0;
    end else begin
      reg_mstatus_spp <= _GEN_320[0];
    end
    if (metaReset) begin
      reg_mstatus_mpie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else if (csr_wen) begin
      if (_T_555) begin
        reg_mstatus_mpie <= _T_3628[7];
      end else if (insn_ret) begin
        if (~io_rw_addr[9]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (!(delegate)) begin
                reg_mstatus_mpie <= reg_mstatus_mie;
              end
            end
          end
        end else if (io_rw_addr[10]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (!(delegate)) begin
                reg_mstatus_mpie <= reg_mstatus_mie;
              end
            end
          end
        end else begin
          reg_mstatus_mpie <= 1'h1;
        end
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (!(delegate)) begin
            reg_mstatus_mpie <= reg_mstatus_mie;
          end
        end
      end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        if (exception) begin
          if (!(trapToDebug)) begin
            if (!(delegate)) begin
              reg_mstatus_mpie <= reg_mstatus_mie;
            end
          end
        end
      end else if (io_rw_addr[10]) begin
        reg_mstatus_mpie <= _GEN_90;
      end else begin
        reg_mstatus_mpie <= 1'h1;
      end
    end else begin
      reg_mstatus_mpie <= _GEN_90;
    end
    if (metaReset) begin
      reg_mstatus_spie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_spie <= 1'h0;
    end else if (csr_wen) begin
      if (_T_662) begin
        reg_mstatus_spie <= _T_3628[5];
      end else if (_T_555) begin
        reg_mstatus_spie <= _T_3628[5];
      end else if (insn_ret) begin
        reg_mstatus_spie <= _GEN_100;
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (delegate) begin
            reg_mstatus_spie <= reg_mstatus_sie;
          end
        end
      end
    end else if (insn_ret) begin
      reg_mstatus_spie <= _GEN_100;
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (delegate) begin
          reg_mstatus_spie <= reg_mstatus_sie;
        end
      end
    end
    if (metaReset) begin
      reg_mstatus_mie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else if (csr_wen) begin
      if (_T_555) begin
        reg_mstatus_mie <= _T_3628[3];
      end else if (insn_ret) begin
        if (~io_rw_addr[9]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              reg_mstatus_mie <= _GEN_56;
            end
          end
        end else if (io_rw_addr[10]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              reg_mstatus_mie <= _GEN_56;
            end
          end
        end else begin
          reg_mstatus_mie <= reg_mstatus_mpie;
        end
      end else if (exception) begin
        if (!(trapToDebug)) begin
          reg_mstatus_mie <= _GEN_56;
        end
      end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        if (exception) begin
          if (!(trapToDebug)) begin
            reg_mstatus_mie <= _GEN_56;
          end
        end
      end else if (io_rw_addr[10]) begin
        reg_mstatus_mie <= _GEN_92;
      end else begin
        reg_mstatus_mie <= reg_mstatus_mpie;
      end
    end else begin
      reg_mstatus_mie <= _GEN_92;
    end
    if (metaReset) begin
      reg_mstatus_sie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_sie <= 1'h0;
    end else if (csr_wen) begin
      if (_T_662) begin
        reg_mstatus_sie <= _T_3628[1];
      end else if (_T_555) begin
        reg_mstatus_sie <= _T_3628[1];
      end else if (insn_ret) begin
        if (~io_rw_addr[9]) begin
          reg_mstatus_sie <= reg_mstatus_spie;
        end else if (exception) begin
          if (!(trapToDebug)) begin
            if (delegate) begin
              reg_mstatus_sie <= 1'h0;
            end
          end
        end
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (delegate) begin
            reg_mstatus_sie <= 1'h0;
          end
        end
      end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        reg_mstatus_sie <= reg_mstatus_spie;
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (delegate) begin
            reg_mstatus_sie <= 1'h0;
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (delegate) begin
          reg_mstatus_sie <= 1'h0;
        end
      end
    end
    if (metaReset) begin
      reg_dcsr_prv <= 2'h0;
    end else if (reset) begin
      reg_dcsr_prv <= 2'h3;
    end else if (csr_wen) begin
      if (_T_564) begin
        if (_T_3748) begin
          reg_dcsr_prv <= 2'h0;
        end else begin
          reg_dcsr_prv <= wdata[1:0];
        end
      end else if (exception) begin
        if (trapToDebug) begin
          if (~reg_debug) begin
            reg_dcsr_prv <= reg_mstatus_prv;
          end
        end
      end
    end else if (exception) begin
      if (trapToDebug) begin
        if (~reg_debug) begin
          reg_dcsr_prv <= reg_mstatus_prv;
        end
      end
    end
    if (metaReset) begin
      reg_singleStepped <= 1'h0;
    end else if (~io_singleStep) begin
      reg_singleStepped <= 1'h0;
    end else begin
      reg_singleStepped <= _GEN_36;
    end
    if (metaReset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else if (reset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else if (csr_wen) begin
      if (_T_564) begin
        reg_dcsr_ebreakm <= wdata[15];
      end
    end
    if (metaReset) begin
      reg_dcsr_ebreaks <= 1'h0;
    end else if (reset) begin
      reg_dcsr_ebreaks <= 1'h0;
    end else if (csr_wen) begin
      if (_T_564) begin
        reg_dcsr_ebreaks <= wdata[13];
      end
    end
    if (metaReset) begin
      reg_dcsr_ebreaku <= 1'h0;
    end else if (reset) begin
      reg_dcsr_ebreaku <= 1'h0;
    end else if (csr_wen) begin
      if (_T_564) begin
        reg_dcsr_ebreaku <= wdata[12];
      end
    end
    if (metaReset) begin
      reg_debug <= 1'h0;
    end else if (reset) begin
      reg_debug <= 1'h0;
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        if (exception) begin
          if (trapToDebug) begin
            reg_debug <= _GEN_38;
          end
        end
      end else if (io_rw_addr[10]) begin
        reg_debug <= 1'h0;
      end else if (exception) begin
        if (trapToDebug) begin
          reg_debug <= _GEN_38;
        end
      end
    end else if (exception) begin
      if (trapToDebug) begin
        reg_debug <= _GEN_38;
      end
    end
    if (metaReset) begin
      reg_mideleg <= 64'h0;
    end else if (csr_wen) begin
      if (_T_672) begin
        reg_mideleg <= wdata;
      end
    end
    if (metaReset) begin
      reg_medeleg <= 64'h0;
    end else if (csr_wen) begin
      if (_T_673) begin
        reg_medeleg <= wdata;
      end
    end
    if (metaReset) begin
      reg_dcsr_cause <= 3'h0;
    end else if (reset) begin
      reg_dcsr_cause <= 3'h0;
    end else if (exception) begin
      if (trapToDebug) begin
        if (~reg_debug) begin
          if (reg_singleStepped) begin
            reg_dcsr_cause <= 3'h4;
          end else begin
            reg_dcsr_cause <= {{1'd0}, _T_1234};
          end
        end
      end
    end
    if (metaReset) begin
      reg_dcsr_step <= 1'h0;
    end else if (reset) begin
      reg_dcsr_step <= 1'h0;
    end else if (csr_wen) begin
      if (_T_564) begin
        reg_dcsr_step <= wdata[2];
      end
    end
    if (metaReset) begin
      reg_dpc <= 40'h0;
    end else begin
      reg_dpc <= _GEN_352[39:0];
    end
    if (metaReset) begin
      reg_dscratch <= 64'h0;
    end else if (csr_wen) begin
      if (_T_566) begin
        reg_dscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_bp_0_control_dmode <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_dmode <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3832) begin
        if (_T_552) begin
          reg_bp_0_control_dmode <= _T_3890;
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_action <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_action <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3832) begin
        if (_T_552) begin
          reg_bp_0_control_action <= _GEN_187;
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_tmatch <= 2'h0;
    end else if (csr_wen) begin
      if (_T_3832) begin
        if (_T_552) begin
          reg_bp_0_control_tmatch <= wdata[8:7];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_m <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3832) begin
        if (_T_552) begin
          reg_bp_0_control_m <= wdata[6];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_s <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3832) begin
        if (_T_552) begin
          reg_bp_0_control_s <= wdata[4];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_u <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3832) begin
        if (_T_552) begin
          reg_bp_0_control_u <= wdata[3];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_x <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3832) begin
        if (_T_552) begin
          reg_bp_0_control_x <= wdata[2];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_w <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3832) begin
        if (_T_552) begin
          reg_bp_0_control_w <= wdata[1];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_r <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3832) begin
        if (_T_552) begin
          reg_bp_0_control_r <= wdata[0];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_address <= 39'h0;
    end else begin
      reg_bp_0_address <= _GEN_366[38:0];
    end
    if (metaReset) begin
      reg_pmp_0_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_0_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3975) begin
        reg_pmp_0_cfg_l <= wdata[7];
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_0_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_3975) begin
        reg_pmp_0_cfg_a <= wdata[4:3];
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3975) begin
        reg_pmp_0_cfg_x <= wdata[2];
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3975) begin
        reg_pmp_0_cfg_w <= _T_3985;
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3975) begin
        reg_pmp_0_cfg_r <= wdata[0];
      end
    end
    if (metaReset) begin
      reg_pmp_0_addr <= 30'h0;
    end else begin
      reg_pmp_0_addr <= _GEN_404[29:0];
    end
    if (metaReset) begin
      reg_pmp_1_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_1_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3995) begin
        reg_pmp_1_cfg_l <= wdata[15];
      end
    end
    if (metaReset) begin
      reg_pmp_1_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_1_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_3995) begin
        reg_pmp_1_cfg_a <= wdata[12:11];
      end
    end
    if (metaReset) begin
      reg_pmp_1_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3995) begin
        reg_pmp_1_cfg_x <= wdata[10];
      end
    end
    if (metaReset) begin
      reg_pmp_1_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3995) begin
        reg_pmp_1_cfg_w <= _T_4005;
      end
    end
    if (metaReset) begin
      reg_pmp_1_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3995) begin
        reg_pmp_1_cfg_r <= wdata[8];
      end
    end
    if (metaReset) begin
      reg_pmp_1_addr <= 30'h0;
    end else begin
      reg_pmp_1_addr <= _GEN_411[29:0];
    end
    if (metaReset) begin
      reg_pmp_2_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_2_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4015) begin
        reg_pmp_2_cfg_l <= wdata[23];
      end
    end
    if (metaReset) begin
      reg_pmp_2_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_2_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_4015) begin
        reg_pmp_2_cfg_a <= wdata[20:19];
      end
    end
    if (metaReset) begin
      reg_pmp_2_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4015) begin
        reg_pmp_2_cfg_x <= wdata[18];
      end
    end
    if (metaReset) begin
      reg_pmp_2_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4015) begin
        reg_pmp_2_cfg_w <= _T_4025;
      end
    end
    if (metaReset) begin
      reg_pmp_2_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4015) begin
        reg_pmp_2_cfg_r <= wdata[16];
      end
    end
    if (metaReset) begin
      reg_pmp_2_addr <= 30'h0;
    end else begin
      reg_pmp_2_addr <= _GEN_418[29:0];
    end
    if (metaReset) begin
      reg_pmp_3_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_3_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4035) begin
        reg_pmp_3_cfg_l <= wdata[31];
      end
    end
    if (metaReset) begin
      reg_pmp_3_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_3_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_4035) begin
        reg_pmp_3_cfg_a <= wdata[28:27];
      end
    end
    if (metaReset) begin
      reg_pmp_3_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4035) begin
        reg_pmp_3_cfg_x <= wdata[26];
      end
    end
    if (metaReset) begin
      reg_pmp_3_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4035) begin
        reg_pmp_3_cfg_w <= _T_4045;
      end
    end
    if (metaReset) begin
      reg_pmp_3_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4035) begin
        reg_pmp_3_cfg_r <= wdata[24];
      end
    end
    if (metaReset) begin
      reg_pmp_3_addr <= 30'h0;
    end else begin
      reg_pmp_3_addr <= _GEN_425[29:0];
    end
    if (metaReset) begin
      reg_pmp_4_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_4_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4055) begin
        reg_pmp_4_cfg_l <= wdata[39];
      end
    end
    if (metaReset) begin
      reg_pmp_4_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_4_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_4055) begin
        reg_pmp_4_cfg_a <= wdata[36:35];
      end
    end
    if (metaReset) begin
      reg_pmp_4_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4055) begin
        reg_pmp_4_cfg_x <= wdata[34];
      end
    end
    if (metaReset) begin
      reg_pmp_4_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4055) begin
        reg_pmp_4_cfg_w <= _T_4065;
      end
    end
    if (metaReset) begin
      reg_pmp_4_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4055) begin
        reg_pmp_4_cfg_r <= wdata[32];
      end
    end
    if (metaReset) begin
      reg_pmp_4_addr <= 30'h0;
    end else begin
      reg_pmp_4_addr <= _GEN_432[29:0];
    end
    if (metaReset) begin
      reg_pmp_5_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_5_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4075) begin
        reg_pmp_5_cfg_l <= wdata[47];
      end
    end
    if (metaReset) begin
      reg_pmp_5_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_5_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_4075) begin
        reg_pmp_5_cfg_a <= wdata[44:43];
      end
    end
    if (metaReset) begin
      reg_pmp_5_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4075) begin
        reg_pmp_5_cfg_x <= wdata[42];
      end
    end
    if (metaReset) begin
      reg_pmp_5_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4075) begin
        reg_pmp_5_cfg_w <= _T_4085;
      end
    end
    if (metaReset) begin
      reg_pmp_5_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4075) begin
        reg_pmp_5_cfg_r <= wdata[40];
      end
    end
    if (metaReset) begin
      reg_pmp_5_addr <= 30'h0;
    end else begin
      reg_pmp_5_addr <= _GEN_439[29:0];
    end
    if (metaReset) begin
      reg_pmp_6_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_6_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4095) begin
        reg_pmp_6_cfg_l <= wdata[55];
      end
    end
    if (metaReset) begin
      reg_pmp_6_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_6_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_4095) begin
        reg_pmp_6_cfg_a <= wdata[52:51];
      end
    end
    if (metaReset) begin
      reg_pmp_6_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4095) begin
        reg_pmp_6_cfg_x <= wdata[50];
      end
    end
    if (metaReset) begin
      reg_pmp_6_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4095) begin
        reg_pmp_6_cfg_w <= _T_4105;
      end
    end
    if (metaReset) begin
      reg_pmp_6_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4095) begin
        reg_pmp_6_cfg_r <= wdata[48];
      end
    end
    if (metaReset) begin
      reg_pmp_6_addr <= 30'h0;
    end else begin
      reg_pmp_6_addr <= _GEN_446[29:0];
    end
    if (metaReset) begin
      reg_pmp_7_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_7_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4115) begin
        reg_pmp_7_cfg_l <= wdata[63];
      end
    end
    if (metaReset) begin
      reg_pmp_7_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_7_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_4115) begin
        reg_pmp_7_cfg_a <= wdata[60:59];
      end
    end
    if (metaReset) begin
      reg_pmp_7_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4115) begin
        reg_pmp_7_cfg_x <= wdata[58];
      end
    end
    if (metaReset) begin
      reg_pmp_7_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4115) begin
        reg_pmp_7_cfg_w <= _T_4125;
      end
    end
    if (metaReset) begin
      reg_pmp_7_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4115) begin
        reg_pmp_7_cfg_r <= wdata[56];
      end
    end
    if (metaReset) begin
      reg_pmp_7_addr <= 30'h0;
    end else begin
      reg_pmp_7_addr <= _GEN_453[29:0];
    end
    if (metaReset) begin
      reg_mie <= 64'h0;
    end else if (csr_wen) begin
      if (_T_664) begin
        reg_mie <= _T_3824;
      end else if (_T_558) begin
        reg_mie <= _T_3721;
      end
    end
    if (metaReset) begin
      reg_mip_seip <= 1'h0;
    end else if (csr_wen) begin
      if (_T_557) begin
        reg_mip_seip <= _T_3702[9];
      end
    end
    if (metaReset) begin
      reg_mip_stip <= 1'h0;
    end else if (csr_wen) begin
      if (_T_557) begin
        reg_mip_stip <= _T_3702[5];
      end
    end
    if (metaReset) begin
      reg_mip_ssip <= 1'h0;
    end else if (csr_wen) begin
      if (_T_663) begin
        reg_mip_ssip <= _T_3792[1];
      end else if (_T_557) begin
        reg_mip_ssip <= _T_3702[1];
      end
    end
    if (metaReset) begin
      reg_mepc <= 40'h0;
    end else begin
      reg_mepc <= _GEN_335[39:0];
    end
    if (metaReset) begin
      reg_mcause <= 64'h0;
    end else if (reset) begin
      reg_mcause <= 64'h0;
    end else if (csr_wen) begin
      if (_T_562) begin
        reg_mcause <= _T_3725;
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (!(delegate)) begin
            if (insn_call) begin
              reg_mcause <= {{60'd0}, _T_1143};
            end else if (insn_break) begin
              reg_mcause <= 64'h3;
            end else begin
              reg_mcause <= io_cause;
            end
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (!(delegate)) begin
          if (insn_call) begin
            reg_mcause <= {{60'd0}, _T_1143};
          end else if (insn_break) begin
            reg_mcause <= 64'h3;
          end else begin
            reg_mcause <= io_cause;
          end
        end
      end
    end
    if (metaReset) begin
      reg_mtval <= 40'h0;
    end else if (csr_wen) begin
      if (_T_561) begin
        reg_mtval <= wdata[39:0];
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (!(delegate)) begin
            reg_mtval <= io_tval;
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (!(delegate)) begin
          reg_mtval <= io_tval;
        end
      end
    end
    if (metaReset) begin
      reg_mscratch <= 64'h0;
    end else if (csr_wen) begin
      if (_T_559) begin
        reg_mscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_mtvec <= 32'h0;
    end else if (reset) begin
      reg_mtvec <= 32'h0;
    end else begin
      reg_mtvec <= _GEN_337[31:0];
    end
    if (metaReset) begin
      reg_mcounteren <= 32'h0;
    end else begin
      reg_mcounteren <= _GEN_364[31:0];
    end
    if (metaReset) begin
      reg_scounteren <= 32'h0;
    end else begin
      reg_scounteren <= _GEN_363[31:0];
    end
    if (metaReset) begin
      reg_sepc <= 40'h0;
    end else begin
      reg_sepc <= _GEN_357[39:0];
    end
    if (metaReset) begin
      reg_scause <= 64'h0;
    end else if (csr_wen) begin
      if (_T_666) begin
        reg_scause <= _T_3828;
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (delegate) begin
            if (insn_call) begin
              reg_scause <= {{60'd0}, _T_1143};
            end else if (insn_break) begin
              reg_scause <= 64'h3;
            end else begin
              reg_scause <= io_cause;
            end
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (delegate) begin
          if (insn_call) begin
            reg_scause <= {{60'd0}, _T_1143};
          end else if (insn_break) begin
            reg_scause <= 64'h3;
          end else begin
            reg_scause <= io_cause;
          end
        end
      end
    end
    if (metaReset) begin
      reg_stval <= 40'h0;
    end else if (csr_wen) begin
      if (_T_667) begin
        reg_stval <= wdata[39:0];
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (delegate) begin
            reg_stval <= io_tval;
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (delegate) begin
          reg_stval <= io_tval;
        end
      end
    end
    if (metaReset) begin
      reg_sscratch <= 64'h0;
    end else if (csr_wen) begin
      if (_T_665) begin
        reg_sscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_stvec <= 39'h0;
    end else begin
      reg_stvec <= _GEN_358[38:0];
    end
    if (metaReset) begin
      reg_satp_mode <= 4'h0;
    end else if (csr_wen) begin
      if (_T_668) begin
        if (_T_3818) begin
          reg_satp_mode <= _T_3819;
        end
      end
    end
    if (metaReset) begin
      reg_satp_ppn <= 44'h0;
    end else if (csr_wen) begin
      if (_T_668) begin
        if (_T_3818) begin
          reg_satp_ppn <= {{24'd0}, wdata[19:0]};
        end
      end
    end
    if (metaReset) begin
      reg_fflags <= 5'h0;
    end else begin
      reg_fflags <= _GEN_345[4:0];
    end
    if (metaReset) begin
      reg_frm <= 3'h0;
    end else begin
      reg_frm <= _GEN_346[2:0];
    end
    if (metaReset) begin
      _T_39 <= 6'h0;
    end else if (reset) begin
      _T_39 <= 6'h0;
    end else begin
      _T_39 <= _GEN_342[5:0];
    end
    if (metaReset) begin
      _T_41 <= 58'h0;
    end else if (reset) begin
      _T_41 <= 58'h0;
    end else if (csr_wen) begin
      if (_T_571) begin
        _T_41 <= wdata[63:6];
      end else if (_T_40[6]) begin
        _T_41 <= _T_44;
      end
    end else if (_T_40[6]) begin
      _T_41 <= _T_44;
    end
    if (metaReset) begin
      reg_misa <= 64'h0;
    end else if (reset) begin
      reg_misa <= 64'h800000000094112d;
    end else if (csr_wen) begin
      if (_T_554) begin
        if (_T_3670) begin
          reg_misa <= _T_3679;
        end
      end
    end
    if (metaReset) begin
      reg_custom_0 <= 64'h0;
    end else if (reset) begin
      reg_custom_0 <= 64'h208;
    end else if (csr_wen) begin
      if (_T_692) begin
        reg_custom_0 <= _T_4137;
      end
    end
    if (metaReset) begin
      _T_1196 <= 2'h0;
    end else if (_T_1194) begin
      _T_1196 <= reg_mstatus_mpp;
    end else begin
      _T_1196 <= reg_mstatus_prv;
    end
    if (metaReset) begin
      _T_1579 <= 1'h0;
    end else if (reset) begin
      _T_1579 <= 1'h0;
    end else begin
      _T_1579 <= _GEN_117;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1206) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:674 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n"); // @[CSR.scala 674:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1206) begin
          $fatal; // @[CSR.scala 674:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1228) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CSR.scala:682 assert(!reg_singleStepped || io.retire === UInt(0))\n"); // @[CSR.scala 682:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1228) begin
          $fatal; // @[CSR.scala 682:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    CSRFile_state <= CSRFile_xor0;
    if (!(CSRFile_cov_read_data)) begin
      CSRFile_covSum <= CSRFile_covSum + 1'h1;
    end
    if (metaReset) begin
      CSRFile_metaAssert <= 1'h0;
    end else begin
      CSRFile_metaAssert <= CSRFile_metaAssert | CSRFile_or0;
    end
  end
  always @(posedge io_ungated_clock) begin
    if (metaReset) begin
      reg_wfi <= 1'h0;
    end else if (reset) begin
      reg_wfi <= 1'h0;
    end else if (_T_1214) begin
      reg_wfi <= 1'h0;
    end else begin
      reg_wfi <= _GEN_34;
    end
    if (metaReset) begin
      _T_47 <= 6'h0;
    end else if (reset) begin
      _T_47 <= 6'h0;
    end else begin
      _T_47 <= _GEN_340[5:0];
    end
    if (metaReset) begin
      _T_49 <= 58'h0;
    end else if (reset) begin
      _T_49 <= 58'h0;
    end else if (csr_wen) begin
      if (_T_570) begin
        _T_49 <= wdata[63:6];
      end else if (_T_48[6]) begin
        _T_49 <= _T_52;
      end
    end else if (_T_48[6]) begin
      _T_49 <= _T_52;
    end
  end
  always @(posedge clock) begin
    if(CSRFile_cov_write_en & CSRFile_cov_write_mask) begin
      CSRFile_cov[CSRFile_cov_write_addr] <= CSRFile_cov_write_data; // @[Coverage map for CSRFile]
    end
  end
endmodule
module BreakpointUnit(
  input         io_status_debug,
  input  [1:0]  io_status_prv,
  input         io_bp_0_control_action,
  input  [1:0]  io_bp_0_control_tmatch,
  input         io_bp_0_control_m,
  input         io_bp_0_control_s,
  input         io_bp_0_control_u,
  input         io_bp_0_control_x,
  input         io_bp_0_control_w,
  input         io_bp_0_control_r,
  input  [38:0] io_bp_0_address,
  input  [38:0] io_pc,
  input  [38:0] io_ea,
  output        io_xcpt_if,
  output        io_xcpt_ld,
  output        io_xcpt_st,
  output        io_debug_if,
  output        io_debug_ld,
  output        io_debug_st,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [3:0] _T_3; // @[Cat.scala 29:58]
  wire [3:0] _T_4; // @[Breakpoint.scala 31:68]
  wire  _T_6; // @[Breakpoint.scala 31:50]
  wire  _T_7; // @[Breakpoint.scala 83:16]
  wire  _T_9; // @[Breakpoint.scala 45:8]
  wire  _T_11; // @[Breakpoint.scala 45:20]
  wire  _T_15; // @[Breakpoint.scala 39:73]
  wire  _T_17; // @[Breakpoint.scala 39:73]
  wire  _T_19; // @[Breakpoint.scala 39:73]
  wire [3:0] _T_22; // @[Cat.scala 29:58]
  wire [38:0] _GEN_11; // @[Breakpoint.scala 42:9]
  wire [38:0] _T_23; // @[Breakpoint.scala 42:9]
  wire [38:0] _T_35; // @[Breakpoint.scala 42:33]
  wire  _T_36; // @[Breakpoint.scala 42:19]
  wire  _T_37; // @[Breakpoint.scala 48:8]
  wire  _T_38; // @[Breakpoint.scala 83:32]
  wire  _T_39; // @[Breakpoint.scala 84:16]
  wire  _T_70; // @[Breakpoint.scala 84:32]
  wire  _T_71; // @[Breakpoint.scala 85:16]
  wire  _T_73; // @[Breakpoint.scala 45:8]
  wire  _T_75; // @[Breakpoint.scala 45:20]
  wire [38:0] _T_87; // @[Breakpoint.scala 42:9]
  wire  _T_100; // @[Breakpoint.scala 42:19]
  wire  _T_101; // @[Breakpoint.scala 48:8]
  wire  _T_102; // @[Breakpoint.scala 85:32]
  wire [29:0] BreakpointUnit_covSum;
  assign _T_3 = {io_bp_0_control_m,1'h0,io_bp_0_control_s,io_bp_0_control_u}; // @[Cat.scala 29:58]
  assign _T_4 = _T_3 >> io_status_prv; // @[Breakpoint.scala 31:68]
  assign _T_6 = ~io_status_debug & _T_4[0]; // @[Breakpoint.scala 31:50]
  assign _T_7 = _T_6 & io_bp_0_control_r; // @[Breakpoint.scala 83:16]
  assign _T_9 = io_ea >= io_bp_0_address; // @[Breakpoint.scala 45:8]
  assign _T_11 = _T_9 ^ io_bp_0_control_tmatch[0]; // @[Breakpoint.scala 45:20]
  assign _T_15 = io_bp_0_control_tmatch[0] & io_bp_0_address[0]; // @[Breakpoint.scala 39:73]
  assign _T_17 = _T_15 & io_bp_0_address[1]; // @[Breakpoint.scala 39:73]
  assign _T_19 = _T_17 & io_bp_0_address[2]; // @[Breakpoint.scala 39:73]
  assign _T_22 = {_T_19,_T_17,_T_15,io_bp_0_control_tmatch[0]}; // @[Cat.scala 29:58]
  assign _GEN_11 = {{35'd0}, _T_22}; // @[Breakpoint.scala 42:9]
  assign _T_23 = ~io_ea | _GEN_11; // @[Breakpoint.scala 42:9]
  assign _T_35 = ~io_bp_0_address | _GEN_11; // @[Breakpoint.scala 42:33]
  assign _T_36 = _T_23 == _T_35; // @[Breakpoint.scala 42:19]
  assign _T_37 = io_bp_0_control_tmatch[1] ? _T_11 : _T_36; // @[Breakpoint.scala 48:8]
  assign _T_38 = _T_7 & _T_37; // @[Breakpoint.scala 83:32]
  assign _T_39 = _T_6 & io_bp_0_control_w; // @[Breakpoint.scala 84:16]
  assign _T_70 = _T_39 & _T_37; // @[Breakpoint.scala 84:32]
  assign _T_71 = _T_6 & io_bp_0_control_x; // @[Breakpoint.scala 85:16]
  assign _T_73 = io_pc >= io_bp_0_address; // @[Breakpoint.scala 45:8]
  assign _T_75 = _T_73 ^ io_bp_0_control_tmatch[0]; // @[Breakpoint.scala 45:20]
  assign _T_87 = ~io_pc | _GEN_11; // @[Breakpoint.scala 42:9]
  assign _T_100 = _T_87 == _T_35; // @[Breakpoint.scala 42:19]
  assign _T_101 = io_bp_0_control_tmatch[1] ? _T_75 : _T_100; // @[Breakpoint.scala 48:8]
  assign _T_102 = _T_71 & _T_101; // @[Breakpoint.scala 85:32]
  assign io_xcpt_if = _T_102 & ~io_bp_0_control_action; // @[Breakpoint.scala 74:14 Breakpoint.scala 97:40]
  assign io_xcpt_ld = _T_38 & ~io_bp_0_control_action; // @[Breakpoint.scala 75:14 Breakpoint.scala 95:40]
  assign io_xcpt_st = _T_70 & ~io_bp_0_control_action; // @[Breakpoint.scala 76:14 Breakpoint.scala 96:40]
  assign io_debug_if = _T_102 & io_bp_0_control_action; // @[Breakpoint.scala 77:15 Breakpoint.scala 97:73]
  assign io_debug_ld = _T_38 & io_bp_0_control_action; // @[Breakpoint.scala 78:15 Breakpoint.scala 95:73]
  assign io_debug_st = _T_70 & io_bp_0_control_action; // @[Breakpoint.scala 79:15 Breakpoint.scala 96:73]
  assign BreakpointUnit_covSum = 30'h0;
  assign io_covSum = BreakpointUnit_covSum;
  assign metaAssert = 1'h0;
endmodule
module ALU(
  input         io_dw,
  input  [3:0]  io_fn,
  input  [63:0] io_in2,
  input  [63:0] io_in1,
  output [63:0] io_out,
  output [63:0] io_adder_out,
  output        io_cmp_out,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [63:0] in2_inv; // @[ALU.scala 62:20]
  wire [63:0] in1_xor_in2; // @[ALU.scala 63:28]
  wire [63:0] _T_3; // @[ALU.scala 64:26]
  wire [63:0] _GEN_1; // @[ALU.scala 64:36]
  wire  _T_9; // @[ALU.scala 68:24]
  wire  _T_14; // @[ALU.scala 69:8]
  wire  slt; // @[ALU.scala 68:8]
  wire  _T_18; // @[ALU.scala 70:68]
  wire  _T_19; // @[ALU.scala 70:41]
  wire  _T_23; // @[ALU.scala 77:46]
  wire [31:0] _T_25; // @[Bitwise.scala 72:12]
  wire [31:0] _T_28; // @[ALU.scala 78:24]
  wire  _T_31; // @[ALU.scala 79:33]
  wire [5:0] shamt; // @[Cat.scala 29:58]
  wire [63:0] shin_r; // @[Cat.scala 29:58]
  wire  _T_34; // @[ALU.scala 82:24]
  wire  _T_35; // @[ALU.scala 82:44]
  wire  _T_36; // @[ALU.scala 82:35]
  wire [63:0] _T_40; // @[Bitwise.scala 103:31]
  wire [63:0] _T_42; // @[Bitwise.scala 103:65]
  wire [63:0] _T_44; // @[Bitwise.scala 103:75]
  wire [63:0] _T_45; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [63:0] _T_50; // @[Bitwise.scala 103:31]
  wire [63:0] _T_52; // @[Bitwise.scala 103:65]
  wire [63:0] _T_54; // @[Bitwise.scala 103:75]
  wire [63:0] _T_55; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_3; // @[Bitwise.scala 103:31]
  wire [63:0] _T_60; // @[Bitwise.scala 103:31]
  wire [63:0] _T_62; // @[Bitwise.scala 103:65]
  wire [63:0] _T_64; // @[Bitwise.scala 103:75]
  wire [63:0] _T_65; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_4; // @[Bitwise.scala 103:31]
  wire [63:0] _T_70; // @[Bitwise.scala 103:31]
  wire [63:0] _T_72; // @[Bitwise.scala 103:65]
  wire [63:0] _T_74; // @[Bitwise.scala 103:75]
  wire [63:0] _T_75; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_5; // @[Bitwise.scala 103:31]
  wire [63:0] _T_80; // @[Bitwise.scala 103:31]
  wire [63:0] _T_82; // @[Bitwise.scala 103:65]
  wire [63:0] _T_84; // @[Bitwise.scala 103:75]
  wire [63:0] _T_85; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_6; // @[Bitwise.scala 103:31]
  wire [63:0] _T_90; // @[Bitwise.scala 103:31]
  wire [63:0] _T_92; // @[Bitwise.scala 103:65]
  wire [63:0] _T_94; // @[Bitwise.scala 103:75]
  wire [63:0] _T_95; // @[Bitwise.scala 103:39]
  wire [63:0] shin; // @[ALU.scala 82:17]
  wire  _T_98; // @[ALU.scala 83:35]
  wire [64:0] _T_100; // @[ALU.scala 83:57]
  wire [64:0] _T_101; // @[ALU.scala 83:64]
  wire [63:0] shout_r; // @[ALU.scala 83:73]
  wire [63:0] _T_105; // @[Bitwise.scala 103:31]
  wire [63:0] _T_107; // @[Bitwise.scala 103:65]
  wire [63:0] _T_109; // @[Bitwise.scala 103:75]
  wire [63:0] _T_110; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_7; // @[Bitwise.scala 103:31]
  wire [63:0] _T_115; // @[Bitwise.scala 103:31]
  wire [63:0] _T_117; // @[Bitwise.scala 103:65]
  wire [63:0] _T_119; // @[Bitwise.scala 103:75]
  wire [63:0] _T_120; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_8; // @[Bitwise.scala 103:31]
  wire [63:0] _T_125; // @[Bitwise.scala 103:31]
  wire [63:0] _T_127; // @[Bitwise.scala 103:65]
  wire [63:0] _T_129; // @[Bitwise.scala 103:75]
  wire [63:0] _T_130; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_9; // @[Bitwise.scala 103:31]
  wire [63:0] _T_135; // @[Bitwise.scala 103:31]
  wire [63:0] _T_137; // @[Bitwise.scala 103:65]
  wire [63:0] _T_139; // @[Bitwise.scala 103:75]
  wire [63:0] _T_140; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_10; // @[Bitwise.scala 103:31]
  wire [63:0] _T_145; // @[Bitwise.scala 103:31]
  wire [63:0] _T_147; // @[Bitwise.scala 103:65]
  wire [63:0] _T_149; // @[Bitwise.scala 103:75]
  wire [63:0] _T_150; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_11; // @[Bitwise.scala 103:31]
  wire [63:0] _T_155; // @[Bitwise.scala 103:31]
  wire [63:0] _T_157; // @[Bitwise.scala 103:65]
  wire [63:0] _T_159; // @[Bitwise.scala 103:75]
  wire [63:0] shout_l; // @[Bitwise.scala 103:39]
  wire [63:0] _T_163; // @[ALU.scala 85:18]
  wire  _T_164; // @[ALU.scala 86:25]
  wire [63:0] _T_165; // @[ALU.scala 86:18]
  wire [63:0] shout; // @[ALU.scala 85:74]
  wire  _T_166; // @[ALU.scala 89:25]
  wire  _T_167; // @[ALU.scala 89:45]
  wire  _T_168; // @[ALU.scala 89:36]
  wire [63:0] _T_169; // @[ALU.scala 89:18]
  wire  _T_171; // @[ALU.scala 90:44]
  wire  _T_172; // @[ALU.scala 90:35]
  wire [63:0] _T_173; // @[ALU.scala 90:63]
  wire [63:0] _T_174; // @[ALU.scala 90:18]
  wire [63:0] logic_; // @[ALU.scala 89:78]
  wire  _T_175; // @[ALU.scala 41:30]
  wire  _T_176; // @[ALU.scala 91:35]
  wire [63:0] _GEN_12; // @[ALU.scala 91:43]
  wire [63:0] _T_177; // @[ALU.scala 91:43]
  wire [63:0] shift_logic; // @[ALU.scala 91:51]
  wire  _T_178; // @[ALU.scala 92:23]
  wire  _T_179; // @[ALU.scala 92:43]
  wire  _T_180; // @[ALU.scala 92:34]
  wire [63:0] out; // @[ALU.scala 92:16]
  wire [31:0] _T_184; // @[Bitwise.scala 72:12]
  wire [63:0] _T_186; // @[Cat.scala 29:58]
  wire [29:0] ALU_covSum;
  assign in2_inv = io_fn[3] ? ~io_in2 : io_in2; // @[ALU.scala 62:20]
  assign in1_xor_in2 = io_in1 ^ in2_inv; // @[ALU.scala 63:28]
  assign _T_3 = io_in1 + in2_inv; // @[ALU.scala 64:26]
  assign _GEN_1 = {{63'd0}, io_fn[3]}; // @[ALU.scala 64:36]
  assign _T_9 = io_in1[63] == io_in2[63]; // @[ALU.scala 68:24]
  assign _T_14 = io_fn[1] ? io_in2[63] : io_in1[63]; // @[ALU.scala 69:8]
  assign slt = _T_9 ? io_adder_out[63] : _T_14; // @[ALU.scala 68:8]
  assign _T_18 = in1_xor_in2 == 64'h0; // @[ALU.scala 70:68]
  assign _T_19 = io_fn[3] ? slt : _T_18; // @[ALU.scala 70:41]
  assign _T_23 = io_fn[3] & io_in1[31]; // @[ALU.scala 77:46]
  assign _T_25 = _T_23 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _T_28 = io_dw ? io_in1[63:32] : _T_25; // @[ALU.scala 78:24]
  assign _T_31 = io_in2[5] & io_dw; // @[ALU.scala 79:33]
  assign shamt = {_T_31,io_in2[4:0]}; // @[Cat.scala 29:58]
  assign shin_r = {_T_28,io_in1[31:0]}; // @[Cat.scala 29:58]
  assign _T_34 = io_fn == 4'h5; // @[ALU.scala 82:24]
  assign _T_35 = io_fn == 4'hb; // @[ALU.scala 82:44]
  assign _T_36 = _T_34 | _T_35; // @[ALU.scala 82:35]
  assign _T_40 = {{32'd0}, shin_r[63:32]}; // @[Bitwise.scala 103:31]
  assign _T_42 = {shin_r[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  assign _T_44 = _T_42 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  assign _T_45 = _T_40 | _T_44; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{16'd0}, _T_45[63:16]}; // @[Bitwise.scala 103:31]
  assign _T_50 = _GEN_2 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  assign _T_52 = {_T_45[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  assign _T_54 = _T_52 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  assign _T_55 = _T_50 | _T_54; // @[Bitwise.scala 103:39]
  assign _GEN_3 = {{8'd0}, _T_55[63:8]}; // @[Bitwise.scala 103:31]
  assign _T_60 = _GEN_3 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  assign _T_62 = {_T_55[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_64 = _T_62 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  assign _T_65 = _T_60 | _T_64; // @[Bitwise.scala 103:39]
  assign _GEN_4 = {{4'd0}, _T_65[63:4]}; // @[Bitwise.scala 103:31]
  assign _T_70 = _GEN_4 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  assign _T_72 = {_T_65[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_74 = _T_72 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  assign _T_75 = _T_70 | _T_74; // @[Bitwise.scala 103:39]
  assign _GEN_5 = {{2'd0}, _T_75[63:2]}; // @[Bitwise.scala 103:31]
  assign _T_80 = _GEN_5 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  assign _T_82 = {_T_75[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_84 = _T_82 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  assign _T_85 = _T_80 | _T_84; // @[Bitwise.scala 103:39]
  assign _GEN_6 = {{1'd0}, _T_85[63:1]}; // @[Bitwise.scala 103:31]
  assign _T_90 = _GEN_6 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  assign _T_92 = {_T_85[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_94 = _T_92 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  assign _T_95 = _T_90 | _T_94; // @[Bitwise.scala 103:39]
  assign shin = _T_36 ? shin_r : _T_95; // @[ALU.scala 82:17]
  assign _T_98 = io_fn[3] & shin[63]; // @[ALU.scala 83:35]
  assign _T_100 = {_T_98,shin}; // @[ALU.scala 83:57]
  assign _T_101 = $signed(_T_100) >>> shamt; // @[ALU.scala 83:64]
  assign shout_r = _T_101[63:0]; // @[ALU.scala 83:73]
  assign _T_105 = {{32'd0}, shout_r[63:32]}; // @[Bitwise.scala 103:31]
  assign _T_107 = {shout_r[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  assign _T_109 = _T_107 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  assign _T_110 = _T_105 | _T_109; // @[Bitwise.scala 103:39]
  assign _GEN_7 = {{16'd0}, _T_110[63:16]}; // @[Bitwise.scala 103:31]
  assign _T_115 = _GEN_7 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  assign _T_117 = {_T_110[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  assign _T_119 = _T_117 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  assign _T_120 = _T_115 | _T_119; // @[Bitwise.scala 103:39]
  assign _GEN_8 = {{8'd0}, _T_120[63:8]}; // @[Bitwise.scala 103:31]
  assign _T_125 = _GEN_8 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  assign _T_127 = {_T_120[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_129 = _T_127 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  assign _T_130 = _T_125 | _T_129; // @[Bitwise.scala 103:39]
  assign _GEN_9 = {{4'd0}, _T_130[63:4]}; // @[Bitwise.scala 103:31]
  assign _T_135 = _GEN_9 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  assign _T_137 = {_T_130[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_139 = _T_137 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  assign _T_140 = _T_135 | _T_139; // @[Bitwise.scala 103:39]
  assign _GEN_10 = {{2'd0}, _T_140[63:2]}; // @[Bitwise.scala 103:31]
  assign _T_145 = _GEN_10 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  assign _T_147 = {_T_140[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_149 = _T_147 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  assign _T_150 = _T_145 | _T_149; // @[Bitwise.scala 103:39]
  assign _GEN_11 = {{1'd0}, _T_150[63:1]}; // @[Bitwise.scala 103:31]
  assign _T_155 = _GEN_11 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  assign _T_157 = {_T_150[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_159 = _T_157 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  assign shout_l = _T_155 | _T_159; // @[Bitwise.scala 103:39]
  assign _T_163 = _T_36 ? shout_r : 64'h0; // @[ALU.scala 85:18]
  assign _T_164 = io_fn == 4'h1; // @[ALU.scala 86:25]
  assign _T_165 = _T_164 ? shout_l : 64'h0; // @[ALU.scala 86:18]
  assign shout = _T_163 | _T_165; // @[ALU.scala 85:74]
  assign _T_166 = io_fn == 4'h4; // @[ALU.scala 89:25]
  assign _T_167 = io_fn == 4'h6; // @[ALU.scala 89:45]
  assign _T_168 = _T_166 | _T_167; // @[ALU.scala 89:36]
  assign _T_169 = _T_168 ? in1_xor_in2 : 64'h0; // @[ALU.scala 89:18]
  assign _T_171 = io_fn == 4'h7; // @[ALU.scala 90:44]
  assign _T_172 = _T_167 | _T_171; // @[ALU.scala 90:35]
  assign _T_173 = io_in1 & io_in2; // @[ALU.scala 90:63]
  assign _T_174 = _T_172 ? _T_173 : 64'h0; // @[ALU.scala 90:18]
  assign logic_ = _T_169 | _T_174; // @[ALU.scala 89:78]
  assign _T_175 = io_fn >= 4'hc; // @[ALU.scala 41:30]
  assign _T_176 = _T_175 & slt; // @[ALU.scala 91:35]
  assign _GEN_12 = {{63'd0}, _T_176}; // @[ALU.scala 91:43]
  assign _T_177 = _GEN_12 | logic_; // @[ALU.scala 91:43]
  assign shift_logic = _T_177 | shout; // @[ALU.scala 91:51]
  assign _T_178 = io_fn == 4'h0; // @[ALU.scala 92:23]
  assign _T_179 = io_fn == 4'ha; // @[ALU.scala 92:43]
  assign _T_180 = _T_178 | _T_179; // @[ALU.scala 92:34]
  assign out = _T_180 ? io_adder_out : shift_logic; // @[ALU.scala 92:16]
  assign _T_184 = out[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _T_186 = {_T_184,out[31:0]}; // @[Cat.scala 29:58]
  assign io_out = io_dw ? out : _T_186; // @[ALU.scala 94:10 ALU.scala 97:37]
  assign io_adder_out = _T_3 + _GEN_1; // @[ALU.scala 64:16]
  assign io_cmp_out = io_fn[0] ^ _T_19; // @[ALU.scala 70:14]
  assign ALU_covSum = 30'h0;
  assign io_covSum = ALU_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulDiv(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [3:0]  io_req_bits_fn,
  input         io_req_bits_dw,
  input  [63:0] io_req_bits_in1,
  input  [63:0] io_req_bits_in2,
  input  [4:0]  io_req_bits_tag,
  input         io_kill,
  input         io_resp_ready,
  output        io_resp_valid,
  output [63:0] io_resp_bits_data,
  output [4:0]  io_resp_bits_tag,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [2:0] state; // @[Multiplier.scala 52:22]
  reg [31:0] _RAND_0;
  reg  req_dw; // @[Multiplier.scala 54:16]
  reg [31:0] _RAND_1;
  reg [4:0] req_tag; // @[Multiplier.scala 54:16]
  reg [31:0] _RAND_2;
  reg [6:0] count; // @[Multiplier.scala 55:18]
  reg [31:0] _RAND_3;
  reg  neg_out; // @[Multiplier.scala 58:20]
  reg [31:0] _RAND_4;
  reg  isHi; // @[Multiplier.scala 59:17]
  reg [31:0] _RAND_5;
  reg  resHi; // @[Multiplier.scala 60:18]
  reg [31:0] _RAND_6;
  reg [64:0] divisor; // @[Multiplier.scala 61:20]
  reg [95:0] _RAND_7;
  reg [129:0] remainder; // @[Multiplier.scala 62:22]
  reg [159:0] _RAND_8;
  wire [3:0] _T; // @[Decode.scala 14:65]
  wire  cmdMul; // @[Decode.scala 14:121]
  wire [3:0] _T_3; // @[Decode.scala 14:65]
  wire  _T_4; // @[Decode.scala 14:121]
  wire [3:0] _T_5; // @[Decode.scala 14:65]
  wire  _T_6; // @[Decode.scala 14:121]
  wire  cmdHi; // @[Decode.scala 15:30]
  wire [3:0] _T_9; // @[Decode.scala 14:65]
  wire  _T_10; // @[Decode.scala 14:121]
  wire [3:0] _T_11; // @[Decode.scala 14:65]
  wire  _T_12; // @[Decode.scala 14:121]
  wire  lhsSigned; // @[Decode.scala 15:30]
  wire  _T_16; // @[Decode.scala 14:121]
  wire  rhsSigned; // @[Decode.scala 15:30]
  wire  _T_23; // @[Multiplier.scala 82:29]
  wire  lhs_sign; // @[Multiplier.scala 82:23]
  wire [31:0] _T_25; // @[Bitwise.scala 72:12]
  wire [31:0] _T_27; // @[Multiplier.scala 83:17]
  wire [63:0] lhs_in; // @[Cat.scala 29:58]
  wire  _T_33; // @[Multiplier.scala 82:29]
  wire  rhs_sign; // @[Multiplier.scala 82:23]
  wire [31:0] _T_35; // @[Bitwise.scala 72:12]
  wire [31:0] _T_37; // @[Multiplier.scala 83:17]
  wire [64:0] subtractor; // @[Multiplier.scala 89:37]
  wire [63:0] result; // @[Multiplier.scala 90:19]
  wire [63:0] negated_remainder; // @[Multiplier.scala 91:27]
  wire  _T_44; // @[Multiplier.scala 93:39]
  wire  _T_47; // @[Multiplier.scala 102:39]
  wire  _T_48; // @[Multiplier.scala 107:39]
  wire [128:0] _T_51; // @[Cat.scala 29:58]
  wire [64:0] _T_55; // @[Multiplier.scala 111:37]
  wire [8:0] _T_59; // @[Multiplier.scala 113:60]
  wire [64:0] _GEN_37; // @[Multiplier.scala 113:67]
  wire [73:0] _T_60; // @[Multiplier.scala 113:67]
  wire [73:0] _GEN_38; // @[Multiplier.scala 113:76]
  wire [73:0] _T_65; // @[Cat.scala 29:58]
  wire [129:0] _T_66; // @[Cat.scala 29:58]
  wire  _T_67; // @[Multiplier.scala 115:32]
  wire  _T_68; // @[Multiplier.scala 115:57]
  wire [10:0] _T_69; // @[Multiplier.scala 117:54]
  wire [64:0] _T_71; // @[Multiplier.scala 117:44]
  wire  _T_73; // @[Multiplier.scala 118:45]
  wire  _T_75; // @[Multiplier.scala 118:79]
  wire  _T_76; // @[Multiplier.scala 118:70]
  wire  _T_78; // @[Multiplier.scala 118:85]
  wire [63:0] _T_80; // @[Multiplier.scala 119:24]
  wire  _T_81; // @[Multiplier.scala 119:37]
  wire  _T_82; // @[Multiplier.scala 119:13]
  wire [10:0] _T_85; // @[Multiplier.scala 120:36]
  wire [128:0] _T_87; // @[Multiplier.scala 120:27]
  wire [129:0] _T_89; // @[Multiplier.scala 121:55]
  wire [128:0] _T_91; // @[Cat.scala 29:58]
  wire [129:0] _T_95; // @[Cat.scala 29:58]
  wire [6:0] _T_97; // @[Multiplier.scala 124:20]
  wire  _T_98; // @[Multiplier.scala 125:25]
  wire  _T_99; // @[Multiplier.scala 125:16]
  wire  _T_100; // @[Multiplier.scala 130:39]
  wire [63:0] _T_104; // @[Multiplier.scala 135:14]
  wire [128:0] _T_108; // @[Cat.scala 29:58]
  wire  _T_109; // @[Multiplier.scala 139:17]
  wire  _T_113; // @[Multiplier.scala 147:24]
  wire  _T_116; // @[Multiplier.scala 147:30]
  wire  _T_121; // @[CircuitMath.scala 37:22]
  wire  _T_124; // @[CircuitMath.scala 37:22]
  wire  _T_127; // @[CircuitMath.scala 37:22]
  wire  _T_130; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_134; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_135; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_139; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_140; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_141; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_142; // @[Cat.scala 29:58]
  wire  _T_145; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_149; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_150; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_154; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_155; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_156; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_157; // @[Cat.scala 29:58]
  wire [2:0] _T_158; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_159; // @[Cat.scala 29:58]
  wire  _T_162; // @[CircuitMath.scala 37:22]
  wire  _T_165; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_169; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_170; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_174; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_175; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_176; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_177; // @[Cat.scala 29:58]
  wire  _T_180; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_184; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_185; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_189; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_190; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_191; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_192; // @[Cat.scala 29:58]
  wire [2:0] _T_193; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_194; // @[Cat.scala 29:58]
  wire [3:0] _T_195; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_196; // @[Cat.scala 29:58]
  wire  _T_199; // @[CircuitMath.scala 37:22]
  wire  _T_202; // @[CircuitMath.scala 37:22]
  wire  _T_205; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_209; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_210; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_214; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_215; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_216; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_217; // @[Cat.scala 29:58]
  wire  _T_220; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_224; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_225; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_229; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_230; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_231; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_232; // @[Cat.scala 29:58]
  wire [2:0] _T_233; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_234; // @[Cat.scala 29:58]
  wire  _T_237; // @[CircuitMath.scala 37:22]
  wire  _T_240; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_244; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_245; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_249; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_250; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_251; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_252; // @[Cat.scala 29:58]
  wire  _T_255; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_259; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_260; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_264; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_265; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_266; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_267; // @[Cat.scala 29:58]
  wire [2:0] _T_268; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_269; // @[Cat.scala 29:58]
  wire [3:0] _T_270; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_271; // @[Cat.scala 29:58]
  wire [4:0] _T_272; // @[CircuitMath.scala 38:21]
  wire [5:0] _T_273; // @[Cat.scala 29:58]
  wire  _T_278; // @[CircuitMath.scala 37:22]
  wire  _T_281; // @[CircuitMath.scala 37:22]
  wire  _T_284; // @[CircuitMath.scala 37:22]
  wire  _T_287; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_291; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_292; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_296; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_297; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_298; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_299; // @[Cat.scala 29:58]
  wire  _T_302; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_306; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_307; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_311; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_312; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_313; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_314; // @[Cat.scala 29:58]
  wire [2:0] _T_315; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_316; // @[Cat.scala 29:58]
  wire  _T_319; // @[CircuitMath.scala 37:22]
  wire  _T_322; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_326; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_327; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_331; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_332; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_333; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_334; // @[Cat.scala 29:58]
  wire  _T_337; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_341; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_342; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_346; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_347; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_348; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_349; // @[Cat.scala 29:58]
  wire [2:0] _T_350; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_351; // @[Cat.scala 29:58]
  wire [3:0] _T_352; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_353; // @[Cat.scala 29:58]
  wire  _T_356; // @[CircuitMath.scala 37:22]
  wire  _T_359; // @[CircuitMath.scala 37:22]
  wire  _T_362; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_366; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_367; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_371; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_372; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_373; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_374; // @[Cat.scala 29:58]
  wire  _T_377; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_381; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_382; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_386; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_387; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_388; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_389; // @[Cat.scala 29:58]
  wire [2:0] _T_390; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_391; // @[Cat.scala 29:58]
  wire  _T_394; // @[CircuitMath.scala 37:22]
  wire  _T_397; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_401; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_402; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_406; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_407; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_408; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_409; // @[Cat.scala 29:58]
  wire  _T_412; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_416; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_417; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_421; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_422; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_423; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_424; // @[Cat.scala 29:58]
  wire [2:0] _T_425; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_426; // @[Cat.scala 29:58]
  wire [3:0] _T_427; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_428; // @[Cat.scala 29:58]
  wire [4:0] _T_429; // @[CircuitMath.scala 38:21]
  wire [5:0] _T_430; // @[Cat.scala 29:58]
  wire [5:0] _T_434; // @[Multiplier.scala 153:35]
  wire  _T_438; // @[Multiplier.scala 154:30]
  wire  _T_439; // @[Multiplier.scala 154:52]
  wire  _T_440; // @[Multiplier.scala 154:41]
  wire [126:0] _GEN_39; // @[Multiplier.scala 156:39]
  wire [126:0] _T_442; // @[Multiplier.scala 156:39]
  wire [128:0] _GEN_16; // @[Multiplier.scala 155:19]
  wire  _T_445; // @[Multiplier.scala 160:18]
  wire  _T_446; // @[Decoupled.scala 40:37]
  wire  _T_447; // @[Multiplier.scala 162:24]
  wire  _T_448; // @[Decoupled.scala 40:37]
  wire  _T_449; // @[Multiplier.scala 166:46]
  wire  _T_454; // @[Multiplier.scala 169:46]
  wire [2:0] _T_455; // @[Multiplier.scala 169:38]
  wire  _T_456; // @[Multiplier.scala 170:46]
  wire [64:0] _T_458; // @[Cat.scala 29:58]
  wire [2:0] _T_460; // @[Multiplier.scala 176:23]
  wire  outMul; // @[Multiplier.scala 176:52]
  wire  _T_466; // @[Multiplier.scala 177:48]
  wire [31:0] loOut; // @[Multiplier.scala 177:18]
  wire [31:0] _T_473; // @[Bitwise.scala 72:12]
  wire [31:0] hiOut; // @[Multiplier.scala 178:18]
  wire  _T_476; // @[Multiplier.scala 182:27]
  wire  _T_477; // @[Multiplier.scala 182:51]
  reg [19:0] MulDiv_state; // @[Register tracking MulDiv state]
  reg [31:0] _RAND_9;
  reg  MulDiv_cov [0:1048575]; // @[Coverage map for MulDiv]
  reg [31:0] _RAND_10;
  wire  MulDiv_cov_read_data; // @[Coverage map for MulDiv]
  wire [19:0] MulDiv_cov_read_addr; // @[Coverage map for MulDiv]
  wire  MulDiv_cov_write_data; // @[Coverage map for MulDiv]
  wire [19:0] MulDiv_cov_write_addr; // @[Coverage map for MulDiv]
  wire  MulDiv_cov_write_mask; // @[Coverage map for MulDiv]
  wire  MulDiv_cov_write_en; // @[Coverage map for MulDiv]
  reg [29:0] MulDiv_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_11;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire  mux_cond_6;
  wire  mux_cond_7;
  wire  mux_cond_8;
  wire  mux_cond_9;
  wire  mux_cond_10;
  wire  mux_cond_11;
  wire  mux_cond_12;
  wire  mux_cond_13;
  wire  mux_cond_14;
  wire  mux_cond_15;
  wire  mux_cond_16;
  wire  mux_cond_17;
  wire  mux_cond_18;
  wire  mux_cond_19;
  wire  mux_cond_20;
  wire  mux_cond_21;
  wire  mux_cond_22;
  wire  mux_cond_23;
  wire  mux_cond_24;
  wire  mux_cond_25;
  wire  mux_cond_26;
  wire  mux_cond_27;
  wire  mux_cond_28;
  wire  mux_cond_29;
  wire  mux_cond_30;
  wire  mux_cond_31;
  wire  mux_cond_32;
  wire  mux_cond_33;
  wire  mux_cond_34;
  wire  mux_cond_35;
  wire  mux_cond_36;
  wire  mux_cond_37;
  wire  mux_cond_38;
  wire  mux_cond_39;
  wire  mux_cond_40;
  wire  mux_cond_41;
  wire  mux_cond_42;
  wire  mux_cond_43;
  wire  mux_cond_44;
  wire  mux_cond_45;
  wire  mux_cond_46;
  wire  mux_cond_47;
  wire  mux_cond_48;
  wire  mux_cond_49;
  wire  mux_cond_50;
  wire  mux_cond_51;
  wire  mux_cond_52;
  wire  mux_cond_53;
  wire  mux_cond_54;
  wire  mux_cond_55;
  wire  mux_cond_56;
  wire  mux_cond_57;
  wire  mux_cond_58;
  wire  mux_cond_59;
  wire  mux_cond_60;
  wire  mux_cond_61;
  wire  mux_cond_62;
  wire  mux_cond_63;
  wire  mux_cond_64;
  wire  mux_cond_65;
  wire  mux_cond_66;
  wire  mux_cond_67;
  wire  mux_cond_68;
  wire  mux_cond_69;
  wire  mux_cond_70;
  wire  mux_cond_71;
  wire  mux_cond_72;
  wire  mux_cond_73;
  wire  mux_cond_74;
  wire  mux_cond_75;
  wire  mux_cond_76;
  wire  mux_cond_77;
  wire  mux_cond_78;
  wire  mux_cond_79;
  wire  mux_cond_80;
  wire  mux_cond_81;
  wire  mux_cond_82;
  wire  mux_cond_83;
  wire  mux_cond_84;
  wire  mux_cond_85;
  wire  mux_cond_86;
  wire  mux_cond_87;
  wire  mux_cond_88;
  wire  mux_cond_89;
  wire  mux_cond_90;
  wire  mux_cond_91;
  wire  mux_cond_92;
  wire  mux_cond_93;
  wire  mux_cond_94;
  wire  mux_cond_95;
  wire  mux_cond_96;
  wire  mux_cond_97;
  wire [6:0] isHi_shl;
  wire [19:0] isHi_pad;
  wire [16:0] neg_out_shl;
  wire [19:0] neg_out_pad;
  wire [14:0] req_dw_shl;
  wire [19:0] req_dw_pad;
  wire [17:0] state_shl;
  wire [19:0] state_pad;
  wire [19:0] resHi_shl;
  wire [19:0] resHi_pad;
  wire [17:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [16:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [13:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [19:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [10:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [11:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [18:0] mux_cond_6_shl;
  wire [19:0] mux_cond_6_pad;
  wire [4:0] mux_cond_7_shl;
  wire [19:0] mux_cond_7_pad;
  wire [14:0] mux_cond_8_shl;
  wire [19:0] mux_cond_8_pad;
  wire [4:0] mux_cond_9_shl;
  wire [19:0] mux_cond_9_pad;
  wire [1:0] mux_cond_10_shl;
  wire [19:0] mux_cond_10_pad;
  wire [19:0] mux_cond_11_shl;
  wire [19:0] mux_cond_11_pad;
  wire [10:0] mux_cond_12_shl;
  wire [19:0] mux_cond_12_pad;
  wire [16:0] mux_cond_13_shl;
  wire [19:0] mux_cond_13_pad;
  wire [9:0] mux_cond_14_shl;
  wire [19:0] mux_cond_14_pad;
  wire [14:0] mux_cond_15_shl;
  wire [19:0] mux_cond_15_pad;
  wire [17:0] mux_cond_16_shl;
  wire [19:0] mux_cond_16_pad;
  wire [4:0] mux_cond_17_shl;
  wire [19:0] mux_cond_17_pad;
  wire [3:0] mux_cond_18_shl;
  wire [19:0] mux_cond_18_pad;
  wire [2:0] mux_cond_19_shl;
  wire [19:0] mux_cond_19_pad;
  wire [15:0] mux_cond_20_shl;
  wire [19:0] mux_cond_20_pad;
  wire [7:0] mux_cond_21_shl;
  wire [19:0] mux_cond_21_pad;
  wire [12:0] mux_cond_22_shl;
  wire [19:0] mux_cond_22_pad;
  wire [13:0] mux_cond_23_shl;
  wire [19:0] mux_cond_23_pad;
  wire [9:0] mux_cond_24_shl;
  wire [19:0] mux_cond_24_pad;
  wire [13:0] mux_cond_25_shl;
  wire [19:0] mux_cond_25_pad;
  wire [17:0] mux_cond_26_shl;
  wire [19:0] mux_cond_26_pad;
  wire [11:0] mux_cond_27_shl;
  wire [19:0] mux_cond_27_pad;
  wire [19:0] mux_cond_28_shl;
  wire [19:0] mux_cond_28_pad;
  wire [2:0] mux_cond_29_shl;
  wire [19:0] mux_cond_29_pad;
  wire [13:0] mux_cond_30_shl;
  wire [19:0] mux_cond_30_pad;
  wire [7:0] mux_cond_31_shl;
  wire [19:0] mux_cond_31_pad;
  wire [16:0] mux_cond_32_shl;
  wire [19:0] mux_cond_32_pad;
  wire [19:0] mux_cond_33_shl;
  wire [19:0] mux_cond_33_pad;
  wire [9:0] mux_cond_34_shl;
  wire [19:0] mux_cond_34_pad;
  wire [9:0] mux_cond_35_shl;
  wire [19:0] mux_cond_35_pad;
  wire [11:0] mux_cond_36_shl;
  wire [19:0] mux_cond_36_pad;
  wire [16:0] mux_cond_37_shl;
  wire [19:0] mux_cond_37_pad;
  wire [2:0] mux_cond_38_shl;
  wire [19:0] mux_cond_38_pad;
  wire [8:0] mux_cond_39_shl;
  wire [19:0] mux_cond_39_pad;
  wire [19:0] mux_cond_40_shl;
  wire [19:0] mux_cond_40_pad;
  wire [12:0] mux_cond_41_shl;
  wire [19:0] mux_cond_41_pad;
  wire [1:0] mux_cond_42_shl;
  wire [19:0] mux_cond_42_pad;
  wire [2:0] mux_cond_43_shl;
  wire [19:0] mux_cond_43_pad;
  wire [10:0] mux_cond_44_shl;
  wire [19:0] mux_cond_44_pad;
  wire [14:0] mux_cond_45_shl;
  wire [19:0] mux_cond_45_pad;
  wire [11:0] mux_cond_46_shl;
  wire [19:0] mux_cond_46_pad;
  wire [11:0] mux_cond_47_shl;
  wire [19:0] mux_cond_47_pad;
  wire [11:0] mux_cond_48_shl;
  wire [19:0] mux_cond_48_pad;
  wire [2:0] mux_cond_49_shl;
  wire [19:0] mux_cond_49_pad;
  wire [9:0] mux_cond_50_shl;
  wire [19:0] mux_cond_50_pad;
  wire [8:0] mux_cond_51_shl;
  wire [19:0] mux_cond_51_pad;
  wire [2:0] mux_cond_52_shl;
  wire [19:0] mux_cond_52_pad;
  wire [7:0] mux_cond_53_shl;
  wire [19:0] mux_cond_53_pad;
  wire [18:0] mux_cond_54_shl;
  wire [19:0] mux_cond_54_pad;
  wire  mux_cond_55_shl;
  wire [19:0] mux_cond_55_pad;
  wire [1:0] mux_cond_56_shl;
  wire [19:0] mux_cond_56_pad;
  wire [15:0] mux_cond_57_shl;
  wire [19:0] mux_cond_57_pad;
  wire [11:0] mux_cond_58_shl;
  wire [19:0] mux_cond_58_pad;
  wire [14:0] mux_cond_59_shl;
  wire [19:0] mux_cond_59_pad;
  wire [12:0] mux_cond_60_shl;
  wire [19:0] mux_cond_60_pad;
  wire [14:0] mux_cond_61_shl;
  wire [19:0] mux_cond_61_pad;
  wire [5:0] mux_cond_62_shl;
  wire [19:0] mux_cond_62_pad;
  wire [6:0] mux_cond_63_shl;
  wire [19:0] mux_cond_63_pad;
  wire [11:0] mux_cond_64_shl;
  wire [19:0] mux_cond_64_pad;
  wire [15:0] mux_cond_65_shl;
  wire [19:0] mux_cond_65_pad;
  wire [18:0] mux_cond_66_shl;
  wire [19:0] mux_cond_66_pad;
  wire [9:0] mux_cond_67_shl;
  wire [19:0] mux_cond_67_pad;
  wire [8:0] mux_cond_68_shl;
  wire [19:0] mux_cond_68_pad;
  wire [2:0] mux_cond_69_shl;
  wire [19:0] mux_cond_69_pad;
  wire [11:0] mux_cond_70_shl;
  wire [19:0] mux_cond_70_pad;
  wire [16:0] mux_cond_71_shl;
  wire [19:0] mux_cond_71_pad;
  wire [16:0] mux_cond_72_shl;
  wire [19:0] mux_cond_72_pad;
  wire [3:0] mux_cond_73_shl;
  wire [19:0] mux_cond_73_pad;
  wire [2:0] mux_cond_74_shl;
  wire [19:0] mux_cond_74_pad;
  wire [4:0] mux_cond_75_shl;
  wire [19:0] mux_cond_75_pad;
  wire [2:0] mux_cond_76_shl;
  wire [19:0] mux_cond_76_pad;
  wire  mux_cond_77_shl;
  wire [19:0] mux_cond_77_pad;
  wire [15:0] mux_cond_78_shl;
  wire [19:0] mux_cond_78_pad;
  wire [2:0] mux_cond_79_shl;
  wire [19:0] mux_cond_79_pad;
  wire [3:0] mux_cond_80_shl;
  wire [19:0] mux_cond_80_pad;
  wire [19:0] mux_cond_81_shl;
  wire [19:0] mux_cond_81_pad;
  wire [9:0] mux_cond_82_shl;
  wire [19:0] mux_cond_82_pad;
  wire [2:0] mux_cond_83_shl;
  wire [19:0] mux_cond_83_pad;
  wire [18:0] mux_cond_84_shl;
  wire [19:0] mux_cond_84_pad;
  wire [2:0] mux_cond_85_shl;
  wire [19:0] mux_cond_85_pad;
  wire [11:0] mux_cond_86_shl;
  wire [19:0] mux_cond_86_pad;
  wire [18:0] mux_cond_87_shl;
  wire [19:0] mux_cond_87_pad;
  wire [8:0] mux_cond_88_shl;
  wire [19:0] mux_cond_88_pad;
  wire [13:0] mux_cond_89_shl;
  wire [19:0] mux_cond_89_pad;
  wire [5:0] mux_cond_90_shl;
  wire [19:0] mux_cond_90_pad;
  wire [5:0] mux_cond_91_shl;
  wire [19:0] mux_cond_91_pad;
  wire [4:0] mux_cond_92_shl;
  wire [19:0] mux_cond_92_pad;
  wire [8:0] mux_cond_93_shl;
  wire [19:0] mux_cond_93_pad;
  wire [17:0] mux_cond_94_shl;
  wire [19:0] mux_cond_94_pad;
  wire [17:0] mux_cond_95_shl;
  wire [19:0] mux_cond_95_pad;
  wire [9:0] mux_cond_96_shl;
  wire [19:0] mux_cond_96_pad;
  wire [18:0] mux_cond_97_shl;
  wire [19:0] mux_cond_97_pad;
  wire [19:0] MulDiv_xor64;
  wire [19:0] MulDiv_xor31;
  wire [19:0] MulDiv_xor66;
  wire [19:0] MulDiv_xor32;
  wire [19:0] MulDiv_xor15;
  wire [19:0] MulDiv_xor68;
  wire [19:0] MulDiv_xor33;
  wire [19:0] MulDiv_xor70;
  wire [19:0] MulDiv_xor34;
  wire [19:0] MulDiv_xor16;
  wire [19:0] MulDiv_xor7;
  wire [19:0] MulDiv_xor72;
  wire [19:0] MulDiv_xor35;
  wire [19:0] MulDiv_xor74;
  wire [19:0] MulDiv_xor36;
  wire [19:0] MulDiv_xor17;
  wire [19:0] MulDiv_xor76;
  wire [19:0] MulDiv_xor37;
  wire [19:0] MulDiv_xor77;
  wire [19:0] MulDiv_xor78;
  wire [19:0] MulDiv_xor38;
  wire [19:0] MulDiv_xor18;
  wire [19:0] MulDiv_xor8;
  wire [19:0] MulDiv_xor3;
  wire [19:0] MulDiv_xor80;
  wire [19:0] MulDiv_xor39;
  wire [19:0] MulDiv_xor82;
  wire [19:0] MulDiv_xor40;
  wire [19:0] MulDiv_xor19;
  wire [19:0] MulDiv_xor84;
  wire [19:0] MulDiv_xor41;
  wire [19:0] MulDiv_xor85;
  wire [19:0] MulDiv_xor86;
  wire [19:0] MulDiv_xor42;
  wire [19:0] MulDiv_xor20;
  wire [19:0] MulDiv_xor9;
  wire [19:0] MulDiv_xor88;
  wire [19:0] MulDiv_xor43;
  wire [19:0] MulDiv_xor90;
  wire [19:0] MulDiv_xor44;
  wire [19:0] MulDiv_xor21;
  wire [19:0] MulDiv_xor92;
  wire [19:0] MulDiv_xor45;
  wire [19:0] MulDiv_xor93;
  wire [19:0] MulDiv_xor94;
  wire [19:0] MulDiv_xor46;
  wire [19:0] MulDiv_xor22;
  wire [19:0] MulDiv_xor10;
  wire [19:0] MulDiv_xor4;
  wire [19:0] MulDiv_xor1;
  wire [19:0] MulDiv_xor96;
  wire [19:0] MulDiv_xor47;
  wire [19:0] MulDiv_xor98;
  wire [19:0] MulDiv_xor48;
  wire [19:0] MulDiv_xor23;
  wire [19:0] MulDiv_xor100;
  wire [19:0] MulDiv_xor49;
  wire [19:0] MulDiv_xor101;
  wire [19:0] MulDiv_xor102;
  wire [19:0] MulDiv_xor50;
  wire [19:0] MulDiv_xor24;
  wire [19:0] MulDiv_xor11;
  wire [19:0] MulDiv_xor104;
  wire [19:0] MulDiv_xor51;
  wire [19:0] MulDiv_xor106;
  wire [19:0] MulDiv_xor52;
  wire [19:0] MulDiv_xor25;
  wire [19:0] MulDiv_xor108;
  wire [19:0] MulDiv_xor53;
  wire [19:0] MulDiv_xor109;
  wire [19:0] MulDiv_xor110;
  wire [19:0] MulDiv_xor54;
  wire [19:0] MulDiv_xor26;
  wire [19:0] MulDiv_xor12;
  wire [19:0] MulDiv_xor5;
  wire [19:0] MulDiv_xor112;
  wire [19:0] MulDiv_xor55;
  wire [19:0] MulDiv_xor114;
  wire [19:0] MulDiv_xor56;
  wire [19:0] MulDiv_xor27;
  wire [19:0] MulDiv_xor116;
  wire [19:0] MulDiv_xor57;
  wire [19:0] MulDiv_xor117;
  wire [19:0] MulDiv_xor118;
  wire [19:0] MulDiv_xor58;
  wire [19:0] MulDiv_xor28;
  wire [19:0] MulDiv_xor13;
  wire [19:0] MulDiv_xor120;
  wire [19:0] MulDiv_xor59;
  wire [19:0] MulDiv_xor122;
  wire [19:0] MulDiv_xor60;
  wire [19:0] MulDiv_xor29;
  wire [19:0] MulDiv_xor124;
  wire [19:0] MulDiv_xor61;
  wire [19:0] MulDiv_xor125;
  wire [19:0] MulDiv_xor126;
  wire [19:0] MulDiv_xor62;
  wire [19:0] MulDiv_xor30;
  wire [19:0] MulDiv_xor14;
  wire [19:0] MulDiv_xor6;
  wire [19:0] MulDiv_xor2;
  wire [19:0] MulDiv_xor0;
  assign _T = io_req_bits_fn & 4'h4; // @[Decode.scala 14:65]
  assign cmdMul = _T == 4'h0; // @[Decode.scala 14:121]
  assign _T_3 = io_req_bits_fn & 4'h5; // @[Decode.scala 14:65]
  assign _T_4 = _T_3 == 4'h1; // @[Decode.scala 14:121]
  assign _T_5 = io_req_bits_fn & 4'h2; // @[Decode.scala 14:65]
  assign _T_6 = _T_5 == 4'h2; // @[Decode.scala 14:121]
  assign cmdHi = _T_4 | _T_6; // @[Decode.scala 15:30]
  assign _T_9 = io_req_bits_fn & 4'h6; // @[Decode.scala 14:65]
  assign _T_10 = _T_9 == 4'h0; // @[Decode.scala 14:121]
  assign _T_11 = io_req_bits_fn & 4'h1; // @[Decode.scala 14:65]
  assign _T_12 = _T_11 == 4'h0; // @[Decode.scala 14:121]
  assign lhsSigned = _T_10 | _T_12; // @[Decode.scala 15:30]
  assign _T_16 = _T_3 == 4'h4; // @[Decode.scala 14:121]
  assign rhsSigned = _T_10 | _T_16; // @[Decode.scala 15:30]
  assign _T_23 = io_req_bits_dw ? io_req_bits_in1[63] : io_req_bits_in1[31]; // @[Multiplier.scala 82:29]
  assign lhs_sign = lhsSigned & _T_23; // @[Multiplier.scala 82:23]
  assign _T_25 = lhs_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _T_27 = io_req_bits_dw ? io_req_bits_in1[63:32] : _T_25; // @[Multiplier.scala 83:17]
  assign lhs_in = {_T_27,io_req_bits_in1[31:0]}; // @[Cat.scala 29:58]
  assign _T_33 = io_req_bits_dw ? io_req_bits_in2[63] : io_req_bits_in2[31]; // @[Multiplier.scala 82:29]
  assign rhs_sign = rhsSigned & _T_33; // @[Multiplier.scala 82:23]
  assign _T_35 = rhs_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _T_37 = io_req_bits_dw ? io_req_bits_in2[63:32] : _T_35; // @[Multiplier.scala 83:17]
  assign subtractor = remainder[128:64] - divisor; // @[Multiplier.scala 89:37]
  assign result = resHi ? remainder[128:65] : remainder[63:0]; // @[Multiplier.scala 90:19]
  assign negated_remainder = 64'h0 - result; // @[Multiplier.scala 91:27]
  assign _T_44 = state == 3'h1; // @[Multiplier.scala 93:39]
  assign _T_47 = state == 3'h5; // @[Multiplier.scala 102:39]
  assign _T_48 = state == 3'h2; // @[Multiplier.scala 107:39]
  assign _T_51 = {remainder[129:65],remainder[63:0]}; // @[Cat.scala 29:58]
  assign _T_55 = _T_51[128:64]; // @[Multiplier.scala 111:37]
  assign _T_59 = {remainder[64],_T_51[7:0]}; // @[Multiplier.scala 113:60]
  assign _GEN_37 = {{56{_T_59[8]}},_T_59}; // @[Multiplier.scala 113:67]
  assign _T_60 = $signed(_GEN_37) * $signed(divisor); // @[Multiplier.scala 113:67]
  assign _GEN_38 = {{9{_T_55[64]}},_T_55}; // @[Multiplier.scala 113:76]
  assign _T_65 = $signed(_T_60) + $signed(_GEN_38); // @[Cat.scala 29:58]
  assign _T_66 = {_T_65,_T_51[63:8]}; // @[Cat.scala 29:58]
  assign _T_67 = count == 7'h6; // @[Multiplier.scala 115:32]
  assign _T_68 = _T_67 & neg_out; // @[Multiplier.scala 115:57]
  assign _T_69 = count * 7'h8; // @[Multiplier.scala 117:54]
  assign _T_71 = -65'sh10000000000000000 >>> _T_69[5:0]; // @[Multiplier.scala 117:44]
  assign _T_73 = count != 7'h7; // @[Multiplier.scala 118:45]
  assign _T_75 = count != 7'h0; // @[Multiplier.scala 118:79]
  assign _T_76 = _T_73 & _T_75; // @[Multiplier.scala 118:70]
  assign _T_78 = _T_76 & ~isHi; // @[Multiplier.scala 118:85]
  assign _T_80 = _T_51[63:0] & ~_T_71[63:0]; // @[Multiplier.scala 119:24]
  assign _T_81 = _T_80 == 64'h0; // @[Multiplier.scala 119:37]
  assign _T_82 = _T_78 & _T_81; // @[Multiplier.scala 119:13]
  assign _T_85 = 11'h40 - _T_69; // @[Multiplier.scala 120:36]
  assign _T_87 = _T_51 >> _T_85[5:0]; // @[Multiplier.scala 120:27]
  assign _T_89 = _T_82 ? {{1'd0}, _T_87} : _T_66; // @[Multiplier.scala 121:55]
  assign _T_91 = {_T_66[128:64],_T_89[63:0]}; // @[Cat.scala 29:58]
  assign _T_95 = {_T_91[128:64],_T_68,_T_91[63:0]}; // @[Cat.scala 29:58]
  assign _T_97 = count + 7'h1; // @[Multiplier.scala 124:20]
  assign _T_98 = count == 7'h7; // @[Multiplier.scala 125:25]
  assign _T_99 = _T_82 | _T_98; // @[Multiplier.scala 125:16]
  assign _T_100 = state == 3'h3; // @[Multiplier.scala 130:39]
  assign _T_104 = subtractor[64] ? remainder[127:64] : subtractor[63:0]; // @[Multiplier.scala 135:14]
  assign _T_108 = {_T_104,remainder[63:0],~subtractor[64]}; // @[Cat.scala 29:58]
  assign _T_109 = count == 7'h40; // @[Multiplier.scala 139:17]
  assign _T_113 = count == 7'h0; // @[Multiplier.scala 147:24]
  assign _T_116 = _T_113 & ~subtractor[64]; // @[Multiplier.scala 147:30]
  assign _T_121 = |divisor[63:32]; // @[CircuitMath.scala 37:22]
  assign _T_124 = |divisor[63:48]; // @[CircuitMath.scala 37:22]
  assign _T_127 = |divisor[63:56]; // @[CircuitMath.scala 37:22]
  assign _T_130 = |divisor[63:60]; // @[CircuitMath.scala 37:22]
  assign _T_134 = divisor[62] ? 2'h2 : {{1'd0}, divisor[61]}; // @[CircuitMath.scala 32:10]
  assign _T_135 = divisor[63] ? 2'h3 : _T_134; // @[CircuitMath.scala 32:10]
  assign _T_139 = divisor[58] ? 2'h2 : {{1'd0}, divisor[57]}; // @[CircuitMath.scala 32:10]
  assign _T_140 = divisor[59] ? 2'h3 : _T_139; // @[CircuitMath.scala 32:10]
  assign _T_141 = _T_130 ? _T_135 : _T_140; // @[CircuitMath.scala 38:21]
  assign _T_142 = {_T_130,_T_141}; // @[Cat.scala 29:58]
  assign _T_145 = |divisor[55:52]; // @[CircuitMath.scala 37:22]
  assign _T_149 = divisor[54] ? 2'h2 : {{1'd0}, divisor[53]}; // @[CircuitMath.scala 32:10]
  assign _T_150 = divisor[55] ? 2'h3 : _T_149; // @[CircuitMath.scala 32:10]
  assign _T_154 = divisor[50] ? 2'h2 : {{1'd0}, divisor[49]}; // @[CircuitMath.scala 32:10]
  assign _T_155 = divisor[51] ? 2'h3 : _T_154; // @[CircuitMath.scala 32:10]
  assign _T_156 = _T_145 ? _T_150 : _T_155; // @[CircuitMath.scala 38:21]
  assign _T_157 = {_T_145,_T_156}; // @[Cat.scala 29:58]
  assign _T_158 = _T_127 ? _T_142 : _T_157; // @[CircuitMath.scala 38:21]
  assign _T_159 = {_T_127,_T_158}; // @[Cat.scala 29:58]
  assign _T_162 = |divisor[47:40]; // @[CircuitMath.scala 37:22]
  assign _T_165 = |divisor[47:44]; // @[CircuitMath.scala 37:22]
  assign _T_169 = divisor[46] ? 2'h2 : {{1'd0}, divisor[45]}; // @[CircuitMath.scala 32:10]
  assign _T_170 = divisor[47] ? 2'h3 : _T_169; // @[CircuitMath.scala 32:10]
  assign _T_174 = divisor[42] ? 2'h2 : {{1'd0}, divisor[41]}; // @[CircuitMath.scala 32:10]
  assign _T_175 = divisor[43] ? 2'h3 : _T_174; // @[CircuitMath.scala 32:10]
  assign _T_176 = _T_165 ? _T_170 : _T_175; // @[CircuitMath.scala 38:21]
  assign _T_177 = {_T_165,_T_176}; // @[Cat.scala 29:58]
  assign _T_180 = |divisor[39:36]; // @[CircuitMath.scala 37:22]
  assign _T_184 = divisor[38] ? 2'h2 : {{1'd0}, divisor[37]}; // @[CircuitMath.scala 32:10]
  assign _T_185 = divisor[39] ? 2'h3 : _T_184; // @[CircuitMath.scala 32:10]
  assign _T_189 = divisor[34] ? 2'h2 : {{1'd0}, divisor[33]}; // @[CircuitMath.scala 32:10]
  assign _T_190 = divisor[35] ? 2'h3 : _T_189; // @[CircuitMath.scala 32:10]
  assign _T_191 = _T_180 ? _T_185 : _T_190; // @[CircuitMath.scala 38:21]
  assign _T_192 = {_T_180,_T_191}; // @[Cat.scala 29:58]
  assign _T_193 = _T_162 ? _T_177 : _T_192; // @[CircuitMath.scala 38:21]
  assign _T_194 = {_T_162,_T_193}; // @[Cat.scala 29:58]
  assign _T_195 = _T_124 ? _T_159 : _T_194; // @[CircuitMath.scala 38:21]
  assign _T_196 = {_T_124,_T_195}; // @[Cat.scala 29:58]
  assign _T_199 = |divisor[31:16]; // @[CircuitMath.scala 37:22]
  assign _T_202 = |divisor[31:24]; // @[CircuitMath.scala 37:22]
  assign _T_205 = |divisor[31:28]; // @[CircuitMath.scala 37:22]
  assign _T_209 = divisor[30] ? 2'h2 : {{1'd0}, divisor[29]}; // @[CircuitMath.scala 32:10]
  assign _T_210 = divisor[31] ? 2'h3 : _T_209; // @[CircuitMath.scala 32:10]
  assign _T_214 = divisor[26] ? 2'h2 : {{1'd0}, divisor[25]}; // @[CircuitMath.scala 32:10]
  assign _T_215 = divisor[27] ? 2'h3 : _T_214; // @[CircuitMath.scala 32:10]
  assign _T_216 = _T_205 ? _T_210 : _T_215; // @[CircuitMath.scala 38:21]
  assign _T_217 = {_T_205,_T_216}; // @[Cat.scala 29:58]
  assign _T_220 = |divisor[23:20]; // @[CircuitMath.scala 37:22]
  assign _T_224 = divisor[22] ? 2'h2 : {{1'd0}, divisor[21]}; // @[CircuitMath.scala 32:10]
  assign _T_225 = divisor[23] ? 2'h3 : _T_224; // @[CircuitMath.scala 32:10]
  assign _T_229 = divisor[18] ? 2'h2 : {{1'd0}, divisor[17]}; // @[CircuitMath.scala 32:10]
  assign _T_230 = divisor[19] ? 2'h3 : _T_229; // @[CircuitMath.scala 32:10]
  assign _T_231 = _T_220 ? _T_225 : _T_230; // @[CircuitMath.scala 38:21]
  assign _T_232 = {_T_220,_T_231}; // @[Cat.scala 29:58]
  assign _T_233 = _T_202 ? _T_217 : _T_232; // @[CircuitMath.scala 38:21]
  assign _T_234 = {_T_202,_T_233}; // @[Cat.scala 29:58]
  assign _T_237 = |divisor[15:8]; // @[CircuitMath.scala 37:22]
  assign _T_240 = |divisor[15:12]; // @[CircuitMath.scala 37:22]
  assign _T_244 = divisor[14] ? 2'h2 : {{1'd0}, divisor[13]}; // @[CircuitMath.scala 32:10]
  assign _T_245 = divisor[15] ? 2'h3 : _T_244; // @[CircuitMath.scala 32:10]
  assign _T_249 = divisor[10] ? 2'h2 : {{1'd0}, divisor[9]}; // @[CircuitMath.scala 32:10]
  assign _T_250 = divisor[11] ? 2'h3 : _T_249; // @[CircuitMath.scala 32:10]
  assign _T_251 = _T_240 ? _T_245 : _T_250; // @[CircuitMath.scala 38:21]
  assign _T_252 = {_T_240,_T_251}; // @[Cat.scala 29:58]
  assign _T_255 = |divisor[7:4]; // @[CircuitMath.scala 37:22]
  assign _T_259 = divisor[6] ? 2'h2 : {{1'd0}, divisor[5]}; // @[CircuitMath.scala 32:10]
  assign _T_260 = divisor[7] ? 2'h3 : _T_259; // @[CircuitMath.scala 32:10]
  assign _T_264 = divisor[2] ? 2'h2 : {{1'd0}, divisor[1]}; // @[CircuitMath.scala 32:10]
  assign _T_265 = divisor[3] ? 2'h3 : _T_264; // @[CircuitMath.scala 32:10]
  assign _T_266 = _T_255 ? _T_260 : _T_265; // @[CircuitMath.scala 38:21]
  assign _T_267 = {_T_255,_T_266}; // @[Cat.scala 29:58]
  assign _T_268 = _T_237 ? _T_252 : _T_267; // @[CircuitMath.scala 38:21]
  assign _T_269 = {_T_237,_T_268}; // @[Cat.scala 29:58]
  assign _T_270 = _T_199 ? _T_234 : _T_269; // @[CircuitMath.scala 38:21]
  assign _T_271 = {_T_199,_T_270}; // @[Cat.scala 29:58]
  assign _T_272 = _T_121 ? _T_196 : _T_271; // @[CircuitMath.scala 38:21]
  assign _T_273 = {_T_121,_T_272}; // @[Cat.scala 29:58]
  assign _T_278 = |remainder[63:32]; // @[CircuitMath.scala 37:22]
  assign _T_281 = |remainder[63:48]; // @[CircuitMath.scala 37:22]
  assign _T_284 = |remainder[63:56]; // @[CircuitMath.scala 37:22]
  assign _T_287 = |remainder[63:60]; // @[CircuitMath.scala 37:22]
  assign _T_291 = remainder[62] ? 2'h2 : {{1'd0}, remainder[61]}; // @[CircuitMath.scala 32:10]
  assign _T_292 = remainder[63] ? 2'h3 : _T_291; // @[CircuitMath.scala 32:10]
  assign _T_296 = remainder[58] ? 2'h2 : {{1'd0}, remainder[57]}; // @[CircuitMath.scala 32:10]
  assign _T_297 = remainder[59] ? 2'h3 : _T_296; // @[CircuitMath.scala 32:10]
  assign _T_298 = _T_287 ? _T_292 : _T_297; // @[CircuitMath.scala 38:21]
  assign _T_299 = {_T_287,_T_298}; // @[Cat.scala 29:58]
  assign _T_302 = |remainder[55:52]; // @[CircuitMath.scala 37:22]
  assign _T_306 = remainder[54] ? 2'h2 : {{1'd0}, remainder[53]}; // @[CircuitMath.scala 32:10]
  assign _T_307 = remainder[55] ? 2'h3 : _T_306; // @[CircuitMath.scala 32:10]
  assign _T_311 = remainder[50] ? 2'h2 : {{1'd0}, remainder[49]}; // @[CircuitMath.scala 32:10]
  assign _T_312 = remainder[51] ? 2'h3 : _T_311; // @[CircuitMath.scala 32:10]
  assign _T_313 = _T_302 ? _T_307 : _T_312; // @[CircuitMath.scala 38:21]
  assign _T_314 = {_T_302,_T_313}; // @[Cat.scala 29:58]
  assign _T_315 = _T_284 ? _T_299 : _T_314; // @[CircuitMath.scala 38:21]
  assign _T_316 = {_T_284,_T_315}; // @[Cat.scala 29:58]
  assign _T_319 = |remainder[47:40]; // @[CircuitMath.scala 37:22]
  assign _T_322 = |remainder[47:44]; // @[CircuitMath.scala 37:22]
  assign _T_326 = remainder[46] ? 2'h2 : {{1'd0}, remainder[45]}; // @[CircuitMath.scala 32:10]
  assign _T_327 = remainder[47] ? 2'h3 : _T_326; // @[CircuitMath.scala 32:10]
  assign _T_331 = remainder[42] ? 2'h2 : {{1'd0}, remainder[41]}; // @[CircuitMath.scala 32:10]
  assign _T_332 = remainder[43] ? 2'h3 : _T_331; // @[CircuitMath.scala 32:10]
  assign _T_333 = _T_322 ? _T_327 : _T_332; // @[CircuitMath.scala 38:21]
  assign _T_334 = {_T_322,_T_333}; // @[Cat.scala 29:58]
  assign _T_337 = |remainder[39:36]; // @[CircuitMath.scala 37:22]
  assign _T_341 = remainder[38] ? 2'h2 : {{1'd0}, remainder[37]}; // @[CircuitMath.scala 32:10]
  assign _T_342 = remainder[39] ? 2'h3 : _T_341; // @[CircuitMath.scala 32:10]
  assign _T_346 = remainder[34] ? 2'h2 : {{1'd0}, remainder[33]}; // @[CircuitMath.scala 32:10]
  assign _T_347 = remainder[35] ? 2'h3 : _T_346; // @[CircuitMath.scala 32:10]
  assign _T_348 = _T_337 ? _T_342 : _T_347; // @[CircuitMath.scala 38:21]
  assign _T_349 = {_T_337,_T_348}; // @[Cat.scala 29:58]
  assign _T_350 = _T_319 ? _T_334 : _T_349; // @[CircuitMath.scala 38:21]
  assign _T_351 = {_T_319,_T_350}; // @[Cat.scala 29:58]
  assign _T_352 = _T_281 ? _T_316 : _T_351; // @[CircuitMath.scala 38:21]
  assign _T_353 = {_T_281,_T_352}; // @[Cat.scala 29:58]
  assign _T_356 = |remainder[31:16]; // @[CircuitMath.scala 37:22]
  assign _T_359 = |remainder[31:24]; // @[CircuitMath.scala 37:22]
  assign _T_362 = |remainder[31:28]; // @[CircuitMath.scala 37:22]
  assign _T_366 = remainder[30] ? 2'h2 : {{1'd0}, remainder[29]}; // @[CircuitMath.scala 32:10]
  assign _T_367 = remainder[31] ? 2'h3 : _T_366; // @[CircuitMath.scala 32:10]
  assign _T_371 = remainder[26] ? 2'h2 : {{1'd0}, remainder[25]}; // @[CircuitMath.scala 32:10]
  assign _T_372 = remainder[27] ? 2'h3 : _T_371; // @[CircuitMath.scala 32:10]
  assign _T_373 = _T_362 ? _T_367 : _T_372; // @[CircuitMath.scala 38:21]
  assign _T_374 = {_T_362,_T_373}; // @[Cat.scala 29:58]
  assign _T_377 = |remainder[23:20]; // @[CircuitMath.scala 37:22]
  assign _T_381 = remainder[22] ? 2'h2 : {{1'd0}, remainder[21]}; // @[CircuitMath.scala 32:10]
  assign _T_382 = remainder[23] ? 2'h3 : _T_381; // @[CircuitMath.scala 32:10]
  assign _T_386 = remainder[18] ? 2'h2 : {{1'd0}, remainder[17]}; // @[CircuitMath.scala 32:10]
  assign _T_387 = remainder[19] ? 2'h3 : _T_386; // @[CircuitMath.scala 32:10]
  assign _T_388 = _T_377 ? _T_382 : _T_387; // @[CircuitMath.scala 38:21]
  assign _T_389 = {_T_377,_T_388}; // @[Cat.scala 29:58]
  assign _T_390 = _T_359 ? _T_374 : _T_389; // @[CircuitMath.scala 38:21]
  assign _T_391 = {_T_359,_T_390}; // @[Cat.scala 29:58]
  assign _T_394 = |remainder[15:8]; // @[CircuitMath.scala 37:22]
  assign _T_397 = |remainder[15:12]; // @[CircuitMath.scala 37:22]
  assign _T_401 = remainder[14] ? 2'h2 : {{1'd0}, remainder[13]}; // @[CircuitMath.scala 32:10]
  assign _T_402 = remainder[15] ? 2'h3 : _T_401; // @[CircuitMath.scala 32:10]
  assign _T_406 = remainder[10] ? 2'h2 : {{1'd0}, remainder[9]}; // @[CircuitMath.scala 32:10]
  assign _T_407 = remainder[11] ? 2'h3 : _T_406; // @[CircuitMath.scala 32:10]
  assign _T_408 = _T_397 ? _T_402 : _T_407; // @[CircuitMath.scala 38:21]
  assign _T_409 = {_T_397,_T_408}; // @[Cat.scala 29:58]
  assign _T_412 = |remainder[7:4]; // @[CircuitMath.scala 37:22]
  assign _T_416 = remainder[6] ? 2'h2 : {{1'd0}, remainder[5]}; // @[CircuitMath.scala 32:10]
  assign _T_417 = remainder[7] ? 2'h3 : _T_416; // @[CircuitMath.scala 32:10]
  assign _T_421 = remainder[2] ? 2'h2 : {{1'd0}, remainder[1]}; // @[CircuitMath.scala 32:10]
  assign _T_422 = remainder[3] ? 2'h3 : _T_421; // @[CircuitMath.scala 32:10]
  assign _T_423 = _T_412 ? _T_417 : _T_422; // @[CircuitMath.scala 38:21]
  assign _T_424 = {_T_412,_T_423}; // @[Cat.scala 29:58]
  assign _T_425 = _T_394 ? _T_409 : _T_424; // @[CircuitMath.scala 38:21]
  assign _T_426 = {_T_394,_T_425}; // @[Cat.scala 29:58]
  assign _T_427 = _T_356 ? _T_391 : _T_426; // @[CircuitMath.scala 38:21]
  assign _T_428 = {_T_356,_T_427}; // @[Cat.scala 29:58]
  assign _T_429 = _T_278 ? _T_353 : _T_428; // @[CircuitMath.scala 38:21]
  assign _T_430 = {_T_278,_T_429}; // @[Cat.scala 29:58]
  assign _T_434 = _T_430 - _T_273; // @[Multiplier.scala 153:35]
  assign _T_438 = _T_113 & ~_T_116; // @[Multiplier.scala 154:30]
  assign _T_439 = ~_T_434 >= 6'h1; // @[Multiplier.scala 154:52]
  assign _T_440 = _T_438 & _T_439; // @[Multiplier.scala 154:41]
  assign _GEN_39 = {{63'd0}, remainder[63:0]}; // @[Multiplier.scala 156:39]
  assign _T_442 = _GEN_39 << ~_T_434; // @[Multiplier.scala 156:39]
  assign _GEN_16 = _T_440 ? {{2'd0}, _T_442} : _T_108; // @[Multiplier.scala 155:19]
  assign _T_445 = _T_116 & ~isHi; // @[Multiplier.scala 160:18]
  assign _T_446 = io_resp_ready & io_resp_valid; // @[Decoupled.scala 40:37]
  assign _T_447 = _T_446 | io_kill; // @[Multiplier.scala 162:24]
  assign _T_448 = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37]
  assign _T_449 = lhs_sign | rhs_sign; // @[Multiplier.scala 166:46]
  assign _T_454 = cmdMul & ~io_req_bits_dw; // @[Multiplier.scala 169:46]
  assign _T_455 = _T_454 ? 3'h4 : 3'h0; // @[Multiplier.scala 169:38]
  assign _T_456 = lhs_sign != rhs_sign; // @[Multiplier.scala 170:46]
  assign _T_458 = {rhs_sign,_T_37,io_req_bits_in2[31:0]}; // @[Cat.scala 29:58]
  assign _T_460 = state & 3'h1; // @[Multiplier.scala 176:23]
  assign outMul = _T_460 == 3'h0; // @[Multiplier.scala 176:52]
  assign _T_466 = ~req_dw & outMul; // @[Multiplier.scala 177:48]
  assign loOut = _T_466 ? result[63:32] : result[31:0]; // @[Multiplier.scala 177:18]
  assign _T_473 = loOut[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign hiOut = req_dw ? result[63:32] : _T_473; // @[Multiplier.scala 178:18]
  assign _T_476 = state == 3'h6; // @[Multiplier.scala 182:27]
  assign _T_477 = state == 3'h7; // @[Multiplier.scala 182:51]
  assign io_req_ready = state == 3'h0; // @[Multiplier.scala 183:16]
  assign io_resp_valid = _T_476 | _T_477; // @[Multiplier.scala 182:17]
  assign io_resp_bits_data = {hiOut,loOut}; // @[Multiplier.scala 181:21]
  assign io_resp_bits_tag = req_tag; // @[Multiplier.scala 179:20]
  assign MulDiv_cov_read_addr = MulDiv_state;
  assign MulDiv_cov_read_data = MulDiv_cov[MulDiv_cov_read_addr]; // @[Coverage map for MulDiv]
  assign MulDiv_cov_write_data = 1'h1;
  assign MulDiv_cov_write_addr = MulDiv_state;
  assign MulDiv_cov_write_mask = 1'h1;
  assign MulDiv_cov_write_en = 1'h1;
  assign mux_cond_0 = remainder[7];
  assign mux_cond_1 = _T_130;
  assign mux_cond_2 = divisor[15];
  assign mux_cond_3 = _T_240;
  assign mux_cond_4 = remainder[38];
  assign mux_cond_5 = _T_205;
  assign mux_cond_6 = remainder[46];
  assign mux_cond_7 = remainder[55];
  assign mux_cond_8 = _T_287;
  assign mux_cond_9 = remainder[62];
  assign mux_cond_10 = divisor[30];
  assign mux_cond_11 = _T_220;
  assign mux_cond_12 = _T_124;
  assign mux_cond_13 = remainder[2];
  assign mux_cond_14 = _T_397;
  assign mux_cond_15 = _T_281;
  assign mux_cond_16 = _T_377;
  assign mux_cond_17 = divisor[63];
  assign mux_cond_18 = remainder[26];
  assign mux_cond_19 = remainder[39];
  assign mux_cond_20 = remainder[54];
  assign mux_cond_21 = remainder[15];
  assign mux_cond_22 = remainder[22];
  assign mux_cond_23 = divisor[18];
  assign mux_cond_24 = divisor[23];
  assign mux_cond_25 = remainder[19];
  assign mux_cond_26 = divisor[22];
  assign mux_cond_27 = remainder[6];
  assign mux_cond_28 = _T_165;
  assign mux_cond_29 = _T_319;
  assign mux_cond_30 = _T_180;
  assign mux_cond_31 = remainder[51];
  assign mux_cond_32 = divisor[50];
  assign mux_cond_33 = divisor[6];
  assign mux_cond_34 = divisor[27];
  assign mux_cond_35 = _T_278;
  assign mux_cond_36 = remainder[47];
  assign mux_cond_37 = remainder[27];
  assign mux_cond_38 = remainder[59];
  assign mux_cond_39 = _T_337;
  assign mux_cond_40 = subtractor[64];
  assign mux_cond_41 = _T_162;
  assign mux_cond_42 = remainder[63];
  assign mux_cond_43 = remainder[3];
  assign mux_cond_44 = remainder[31];
  assign mux_cond_45 = divisor[39];
  assign mux_cond_46 = remainder[18];
  assign mux_cond_47 = remainder[11];
  assign mux_cond_48 = divisor[46];
  assign mux_cond_49 = remainder[34];
  assign mux_cond_50 = divisor[3];
  assign mux_cond_51 = divisor[26];
  assign mux_cond_52 = divisor[54];
  assign mux_cond_53 = remainder[35];
  assign mux_cond_54 = _T_255;
  assign mux_cond_55 = divisor[19];
  assign mux_cond_56 = _T_359;
  assign mux_cond_57 = _T_127;
  assign mux_cond_58 = divisor[11];
  assign mux_cond_59 = _T_145;
  assign mux_cond_60 = divisor[47];
  assign mux_cond_61 = divisor[7];
  assign mux_cond_62 = divisor[34];
  assign mux_cond_63 = divisor[43];
  assign mux_cond_64 = divisor[38];
  assign mux_cond_65 = remainder[58];
  assign mux_cond_66 = divisor[62];
  assign mux_cond_67 = remainder[30];
  assign mux_cond_68 = remainder[63];
  assign mux_cond_69 = _T_202;
  assign mux_cond_70 = _T_199;
  assign mux_cond_71 = _T_302;
  assign mux_cond_72 = divisor[31];
  assign mux_cond_73 = _T_362;
  assign mux_cond_74 = divisor[55];
  assign mux_cond_75 = divisor[63];
  assign mux_cond_76 = remainder[50];
  assign mux_cond_77 = _T_322;
  assign mux_cond_78 = divisor[14];
  assign mux_cond_79 = remainder[14];
  assign mux_cond_80 = remainder[23];
  assign mux_cond_81 = divisor[51];
  assign mux_cond_82 = divisor[10];
  assign mux_cond_83 = remainder[10];
  assign mux_cond_84 = remainder[43];
  assign mux_cond_85 = _T_356;
  assign mux_cond_86 = divisor[35];
  assign mux_cond_87 = remainder[42];
  assign mux_cond_88 = divisor[42];
  assign mux_cond_89 = divisor[58];
  assign mux_cond_90 = _T_412;
  assign mux_cond_91 = divisor[59];
  assign mux_cond_92 = _T_394;
  assign mux_cond_93 = divisor[2];
  assign mux_cond_94 = loOut[31];
  assign mux_cond_95 = _T_237;
  assign mux_cond_96 = _T_121;
  assign mux_cond_97 = _T_284;
  assign isHi_shl = {isHi, 6'h0};
  assign isHi_pad = {13'h0,isHi_shl};
  assign neg_out_shl = {neg_out, 16'h0};
  assign neg_out_pad = {3'h0,neg_out_shl};
  assign req_dw_shl = {req_dw, 14'h0};
  assign req_dw_pad = {5'h0,req_dw_shl};
  assign state_shl = {state, 15'h0};
  assign state_pad = {2'h0,state_shl};
  assign resHi_shl = {resHi, 19'h0};
  assign resHi_pad = resHi_shl;
  assign mux_cond_0_shl = {mux_cond_0, 17'h0};
  assign mux_cond_0_pad = {2'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 16'h0};
  assign mux_cond_1_pad = {3'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 13'h0};
  assign mux_cond_2_pad = {6'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 19'h0};
  assign mux_cond_3_pad = mux_cond_3_shl;
  assign mux_cond_4_shl = {mux_cond_4, 10'h0};
  assign mux_cond_4_pad = {9'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 11'h0};
  assign mux_cond_5_pad = {8'h0,mux_cond_5_shl};
  assign mux_cond_6_shl = {mux_cond_6, 18'h0};
  assign mux_cond_6_pad = {1'h0,mux_cond_6_shl};
  assign mux_cond_7_shl = {mux_cond_7, 4'h0};
  assign mux_cond_7_pad = {15'h0,mux_cond_7_shl};
  assign mux_cond_8_shl = {mux_cond_8, 14'h0};
  assign mux_cond_8_pad = {5'h0,mux_cond_8_shl};
  assign mux_cond_9_shl = {mux_cond_9, 4'h0};
  assign mux_cond_9_pad = {15'h0,mux_cond_9_shl};
  assign mux_cond_10_shl = {mux_cond_10, 1'h0};
  assign mux_cond_10_pad = {18'h0,mux_cond_10_shl};
  assign mux_cond_11_shl = {mux_cond_11, 19'h0};
  assign mux_cond_11_pad = mux_cond_11_shl;
  assign mux_cond_12_shl = {mux_cond_12, 10'h0};
  assign mux_cond_12_pad = {9'h0,mux_cond_12_shl};
  assign mux_cond_13_shl = {mux_cond_13, 16'h0};
  assign mux_cond_13_pad = {3'h0,mux_cond_13_shl};
  assign mux_cond_14_shl = {mux_cond_14, 9'h0};
  assign mux_cond_14_pad = {10'h0,mux_cond_14_shl};
  assign mux_cond_15_shl = {mux_cond_15, 14'h0};
  assign mux_cond_15_pad = {5'h0,mux_cond_15_shl};
  assign mux_cond_16_shl = {mux_cond_16, 17'h0};
  assign mux_cond_16_pad = {2'h0,mux_cond_16_shl};
  assign mux_cond_17_shl = {mux_cond_17, 4'h0};
  assign mux_cond_17_pad = {15'h0,mux_cond_17_shl};
  assign mux_cond_18_shl = {mux_cond_18, 3'h0};
  assign mux_cond_18_pad = {16'h0,mux_cond_18_shl};
  assign mux_cond_19_shl = {mux_cond_19, 2'h0};
  assign mux_cond_19_pad = {17'h0,mux_cond_19_shl};
  assign mux_cond_20_shl = {mux_cond_20, 15'h0};
  assign mux_cond_20_pad = {4'h0,mux_cond_20_shl};
  assign mux_cond_21_shl = {mux_cond_21, 7'h0};
  assign mux_cond_21_pad = {12'h0,mux_cond_21_shl};
  assign mux_cond_22_shl = {mux_cond_22, 12'h0};
  assign mux_cond_22_pad = {7'h0,mux_cond_22_shl};
  assign mux_cond_23_shl = {mux_cond_23, 13'h0};
  assign mux_cond_23_pad = {6'h0,mux_cond_23_shl};
  assign mux_cond_24_shl = {mux_cond_24, 9'h0};
  assign mux_cond_24_pad = {10'h0,mux_cond_24_shl};
  assign mux_cond_25_shl = {mux_cond_25, 13'h0};
  assign mux_cond_25_pad = {6'h0,mux_cond_25_shl};
  assign mux_cond_26_shl = {mux_cond_26, 17'h0};
  assign mux_cond_26_pad = {2'h0,mux_cond_26_shl};
  assign mux_cond_27_shl = {mux_cond_27, 11'h0};
  assign mux_cond_27_pad = {8'h0,mux_cond_27_shl};
  assign mux_cond_28_shl = {mux_cond_28, 19'h0};
  assign mux_cond_28_pad = mux_cond_28_shl;
  assign mux_cond_29_shl = {mux_cond_29, 2'h0};
  assign mux_cond_29_pad = {17'h0,mux_cond_29_shl};
  assign mux_cond_30_shl = {mux_cond_30, 13'h0};
  assign mux_cond_30_pad = {6'h0,mux_cond_30_shl};
  assign mux_cond_31_shl = {mux_cond_31, 7'h0};
  assign mux_cond_31_pad = {12'h0,mux_cond_31_shl};
  assign mux_cond_32_shl = {mux_cond_32, 16'h0};
  assign mux_cond_32_pad = {3'h0,mux_cond_32_shl};
  assign mux_cond_33_shl = {mux_cond_33, 19'h0};
  assign mux_cond_33_pad = mux_cond_33_shl;
  assign mux_cond_34_shl = {mux_cond_34, 9'h0};
  assign mux_cond_34_pad = {10'h0,mux_cond_34_shl};
  assign mux_cond_35_shl = {mux_cond_35, 9'h0};
  assign mux_cond_35_pad = {10'h0,mux_cond_35_shl};
  assign mux_cond_36_shl = {mux_cond_36, 11'h0};
  assign mux_cond_36_pad = {8'h0,mux_cond_36_shl};
  assign mux_cond_37_shl = {mux_cond_37, 16'h0};
  assign mux_cond_37_pad = {3'h0,mux_cond_37_shl};
  assign mux_cond_38_shl = {mux_cond_38, 2'h0};
  assign mux_cond_38_pad = {17'h0,mux_cond_38_shl};
  assign mux_cond_39_shl = {mux_cond_39, 8'h0};
  assign mux_cond_39_pad = {11'h0,mux_cond_39_shl};
  assign mux_cond_40_shl = {mux_cond_40, 19'h0};
  assign mux_cond_40_pad = mux_cond_40_shl;
  assign mux_cond_41_shl = {mux_cond_41, 12'h0};
  assign mux_cond_41_pad = {7'h0,mux_cond_41_shl};
  assign mux_cond_42_shl = {mux_cond_42, 1'h0};
  assign mux_cond_42_pad = {18'h0,mux_cond_42_shl};
  assign mux_cond_43_shl = {mux_cond_43, 2'h0};
  assign mux_cond_43_pad = {17'h0,mux_cond_43_shl};
  assign mux_cond_44_shl = {mux_cond_44, 10'h0};
  assign mux_cond_44_pad = {9'h0,mux_cond_44_shl};
  assign mux_cond_45_shl = {mux_cond_45, 14'h0};
  assign mux_cond_45_pad = {5'h0,mux_cond_45_shl};
  assign mux_cond_46_shl = {mux_cond_46, 11'h0};
  assign mux_cond_46_pad = {8'h0,mux_cond_46_shl};
  assign mux_cond_47_shl = {mux_cond_47, 11'h0};
  assign mux_cond_47_pad = {8'h0,mux_cond_47_shl};
  assign mux_cond_48_shl = {mux_cond_48, 11'h0};
  assign mux_cond_48_pad = {8'h0,mux_cond_48_shl};
  assign mux_cond_49_shl = {mux_cond_49, 2'h0};
  assign mux_cond_49_pad = {17'h0,mux_cond_49_shl};
  assign mux_cond_50_shl = {mux_cond_50, 9'h0};
  assign mux_cond_50_pad = {10'h0,mux_cond_50_shl};
  assign mux_cond_51_shl = {mux_cond_51, 8'h0};
  assign mux_cond_51_pad = {11'h0,mux_cond_51_shl};
  assign mux_cond_52_shl = {mux_cond_52, 2'h0};
  assign mux_cond_52_pad = {17'h0,mux_cond_52_shl};
  assign mux_cond_53_shl = {mux_cond_53, 7'h0};
  assign mux_cond_53_pad = {12'h0,mux_cond_53_shl};
  assign mux_cond_54_shl = {mux_cond_54, 18'h0};
  assign mux_cond_54_pad = {1'h0,mux_cond_54_shl};
  assign mux_cond_55_shl = mux_cond_55;
  assign mux_cond_55_pad = {19'h0,mux_cond_55_shl};
  assign mux_cond_56_shl = {mux_cond_56, 1'h0};
  assign mux_cond_56_pad = {18'h0,mux_cond_56_shl};
  assign mux_cond_57_shl = {mux_cond_57, 15'h0};
  assign mux_cond_57_pad = {4'h0,mux_cond_57_shl};
  assign mux_cond_58_shl = {mux_cond_58, 11'h0};
  assign mux_cond_58_pad = {8'h0,mux_cond_58_shl};
  assign mux_cond_59_shl = {mux_cond_59, 14'h0};
  assign mux_cond_59_pad = {5'h0,mux_cond_59_shl};
  assign mux_cond_60_shl = {mux_cond_60, 12'h0};
  assign mux_cond_60_pad = {7'h0,mux_cond_60_shl};
  assign mux_cond_61_shl = {mux_cond_61, 14'h0};
  assign mux_cond_61_pad = {5'h0,mux_cond_61_shl};
  assign mux_cond_62_shl = {mux_cond_62, 5'h0};
  assign mux_cond_62_pad = {14'h0,mux_cond_62_shl};
  assign mux_cond_63_shl = {mux_cond_63, 6'h0};
  assign mux_cond_63_pad = {13'h0,mux_cond_63_shl};
  assign mux_cond_64_shl = {mux_cond_64, 11'h0};
  assign mux_cond_64_pad = {8'h0,mux_cond_64_shl};
  assign mux_cond_65_shl = {mux_cond_65, 15'h0};
  assign mux_cond_65_pad = {4'h0,mux_cond_65_shl};
  assign mux_cond_66_shl = {mux_cond_66, 18'h0};
  assign mux_cond_66_pad = {1'h0,mux_cond_66_shl};
  assign mux_cond_67_shl = {mux_cond_67, 9'h0};
  assign mux_cond_67_pad = {10'h0,mux_cond_67_shl};
  assign mux_cond_68_shl = {mux_cond_68, 8'h0};
  assign mux_cond_68_pad = {11'h0,mux_cond_68_shl};
  assign mux_cond_69_shl = {mux_cond_69, 2'h0};
  assign mux_cond_69_pad = {17'h0,mux_cond_69_shl};
  assign mux_cond_70_shl = {mux_cond_70, 11'h0};
  assign mux_cond_70_pad = {8'h0,mux_cond_70_shl};
  assign mux_cond_71_shl = {mux_cond_71, 16'h0};
  assign mux_cond_71_pad = {3'h0,mux_cond_71_shl};
  assign mux_cond_72_shl = {mux_cond_72, 16'h0};
  assign mux_cond_72_pad = {3'h0,mux_cond_72_shl};
  assign mux_cond_73_shl = {mux_cond_73, 3'h0};
  assign mux_cond_73_pad = {16'h0,mux_cond_73_shl};
  assign mux_cond_74_shl = {mux_cond_74, 2'h0};
  assign mux_cond_74_pad = {17'h0,mux_cond_74_shl};
  assign mux_cond_75_shl = {mux_cond_75, 4'h0};
  assign mux_cond_75_pad = {15'h0,mux_cond_75_shl};
  assign mux_cond_76_shl = {mux_cond_76, 2'h0};
  assign mux_cond_76_pad = {17'h0,mux_cond_76_shl};
  assign mux_cond_77_shl = mux_cond_77;
  assign mux_cond_77_pad = {19'h0,mux_cond_77_shl};
  assign mux_cond_78_shl = {mux_cond_78, 15'h0};
  assign mux_cond_78_pad = {4'h0,mux_cond_78_shl};
  assign mux_cond_79_shl = {mux_cond_79, 2'h0};
  assign mux_cond_79_pad = {17'h0,mux_cond_79_shl};
  assign mux_cond_80_shl = {mux_cond_80, 3'h0};
  assign mux_cond_80_pad = {16'h0,mux_cond_80_shl};
  assign mux_cond_81_shl = {mux_cond_81, 19'h0};
  assign mux_cond_81_pad = mux_cond_81_shl;
  assign mux_cond_82_shl = {mux_cond_82, 9'h0};
  assign mux_cond_82_pad = {10'h0,mux_cond_82_shl};
  assign mux_cond_83_shl = {mux_cond_83, 2'h0};
  assign mux_cond_83_pad = {17'h0,mux_cond_83_shl};
  assign mux_cond_84_shl = {mux_cond_84, 18'h0};
  assign mux_cond_84_pad = {1'h0,mux_cond_84_shl};
  assign mux_cond_85_shl = {mux_cond_85, 2'h0};
  assign mux_cond_85_pad = {17'h0,mux_cond_85_shl};
  assign mux_cond_86_shl = {mux_cond_86, 11'h0};
  assign mux_cond_86_pad = {8'h0,mux_cond_86_shl};
  assign mux_cond_87_shl = {mux_cond_87, 18'h0};
  assign mux_cond_87_pad = {1'h0,mux_cond_87_shl};
  assign mux_cond_88_shl = {mux_cond_88, 8'h0};
  assign mux_cond_88_pad = {11'h0,mux_cond_88_shl};
  assign mux_cond_89_shl = {mux_cond_89, 13'h0};
  assign mux_cond_89_pad = {6'h0,mux_cond_89_shl};
  assign mux_cond_90_shl = {mux_cond_90, 5'h0};
  assign mux_cond_90_pad = {14'h0,mux_cond_90_shl};
  assign mux_cond_91_shl = {mux_cond_91, 5'h0};
  assign mux_cond_91_pad = {14'h0,mux_cond_91_shl};
  assign mux_cond_92_shl = {mux_cond_92, 4'h0};
  assign mux_cond_92_pad = {15'h0,mux_cond_92_shl};
  assign mux_cond_93_shl = {mux_cond_93, 8'h0};
  assign mux_cond_93_pad = {11'h0,mux_cond_93_shl};
  assign mux_cond_94_shl = {mux_cond_94, 17'h0};
  assign mux_cond_94_pad = {2'h0,mux_cond_94_shl};
  assign mux_cond_95_shl = {mux_cond_95, 17'h0};
  assign mux_cond_95_pad = {2'h0,mux_cond_95_shl};
  assign mux_cond_96_shl = {mux_cond_96, 9'h0};
  assign mux_cond_96_pad = {10'h0,mux_cond_96_shl};
  assign mux_cond_97_shl = {mux_cond_97, 18'h0};
  assign mux_cond_97_pad = {1'h0,mux_cond_97_shl};
  assign MulDiv_xor64 = neg_out_pad ^ req_dw_pad;
  assign MulDiv_xor31 = isHi_pad ^ MulDiv_xor64;
  assign MulDiv_xor66 = resHi_pad ^ mux_cond_0_pad;
  assign MulDiv_xor32 = state_pad ^ MulDiv_xor66;
  assign MulDiv_xor15 = MulDiv_xor31 ^ MulDiv_xor32;
  assign MulDiv_xor68 = mux_cond_2_pad ^ mux_cond_3_pad;
  assign MulDiv_xor33 = mux_cond_1_pad ^ MulDiv_xor68;
  assign MulDiv_xor70 = mux_cond_5_pad ^ mux_cond_6_pad;
  assign MulDiv_xor34 = mux_cond_4_pad ^ MulDiv_xor70;
  assign MulDiv_xor16 = MulDiv_xor33 ^ MulDiv_xor34;
  assign MulDiv_xor7 = MulDiv_xor15 ^ MulDiv_xor16;
  assign MulDiv_xor72 = mux_cond_8_pad ^ mux_cond_9_pad;
  assign MulDiv_xor35 = mux_cond_7_pad ^ MulDiv_xor72;
  assign MulDiv_xor74 = mux_cond_11_pad ^ mux_cond_12_pad;
  assign MulDiv_xor36 = mux_cond_10_pad ^ MulDiv_xor74;
  assign MulDiv_xor17 = MulDiv_xor35 ^ MulDiv_xor36;
  assign MulDiv_xor76 = mux_cond_14_pad ^ mux_cond_15_pad;
  assign MulDiv_xor37 = mux_cond_13_pad ^ MulDiv_xor76;
  assign MulDiv_xor77 = mux_cond_16_pad ^ mux_cond_17_pad;
  assign MulDiv_xor78 = mux_cond_18_pad ^ mux_cond_19_pad;
  assign MulDiv_xor38 = MulDiv_xor77 ^ MulDiv_xor78;
  assign MulDiv_xor18 = MulDiv_xor37 ^ MulDiv_xor38;
  assign MulDiv_xor8 = MulDiv_xor17 ^ MulDiv_xor18;
  assign MulDiv_xor3 = MulDiv_xor7 ^ MulDiv_xor8;
  assign MulDiv_xor80 = mux_cond_21_pad ^ mux_cond_22_pad;
  assign MulDiv_xor39 = mux_cond_20_pad ^ MulDiv_xor80;
  assign MulDiv_xor82 = mux_cond_24_pad ^ mux_cond_25_pad;
  assign MulDiv_xor40 = mux_cond_23_pad ^ MulDiv_xor82;
  assign MulDiv_xor19 = MulDiv_xor39 ^ MulDiv_xor40;
  assign MulDiv_xor84 = mux_cond_27_pad ^ mux_cond_28_pad;
  assign MulDiv_xor41 = mux_cond_26_pad ^ MulDiv_xor84;
  assign MulDiv_xor85 = mux_cond_29_pad ^ mux_cond_30_pad;
  assign MulDiv_xor86 = mux_cond_31_pad ^ mux_cond_32_pad;
  assign MulDiv_xor42 = MulDiv_xor85 ^ MulDiv_xor86;
  assign MulDiv_xor20 = MulDiv_xor41 ^ MulDiv_xor42;
  assign MulDiv_xor9 = MulDiv_xor19 ^ MulDiv_xor20;
  assign MulDiv_xor88 = mux_cond_34_pad ^ mux_cond_35_pad;
  assign MulDiv_xor43 = mux_cond_33_pad ^ MulDiv_xor88;
  assign MulDiv_xor90 = mux_cond_37_pad ^ mux_cond_38_pad;
  assign MulDiv_xor44 = mux_cond_36_pad ^ MulDiv_xor90;
  assign MulDiv_xor21 = MulDiv_xor43 ^ MulDiv_xor44;
  assign MulDiv_xor92 = mux_cond_40_pad ^ mux_cond_41_pad;
  assign MulDiv_xor45 = mux_cond_39_pad ^ MulDiv_xor92;
  assign MulDiv_xor93 = mux_cond_42_pad ^ mux_cond_43_pad;
  assign MulDiv_xor94 = mux_cond_44_pad ^ mux_cond_45_pad;
  assign MulDiv_xor46 = MulDiv_xor93 ^ MulDiv_xor94;
  assign MulDiv_xor22 = MulDiv_xor45 ^ MulDiv_xor46;
  assign MulDiv_xor10 = MulDiv_xor21 ^ MulDiv_xor22;
  assign MulDiv_xor4 = MulDiv_xor9 ^ MulDiv_xor10;
  assign MulDiv_xor1 = MulDiv_xor3 ^ MulDiv_xor4;
  assign MulDiv_xor96 = mux_cond_47_pad ^ mux_cond_48_pad;
  assign MulDiv_xor47 = mux_cond_46_pad ^ MulDiv_xor96;
  assign MulDiv_xor98 = mux_cond_50_pad ^ mux_cond_51_pad;
  assign MulDiv_xor48 = mux_cond_49_pad ^ MulDiv_xor98;
  assign MulDiv_xor23 = MulDiv_xor47 ^ MulDiv_xor48;
  assign MulDiv_xor100 = mux_cond_53_pad ^ mux_cond_54_pad;
  assign MulDiv_xor49 = mux_cond_52_pad ^ MulDiv_xor100;
  assign MulDiv_xor101 = mux_cond_55_pad ^ mux_cond_56_pad;
  assign MulDiv_xor102 = mux_cond_57_pad ^ mux_cond_58_pad;
  assign MulDiv_xor50 = MulDiv_xor101 ^ MulDiv_xor102;
  assign MulDiv_xor24 = MulDiv_xor49 ^ MulDiv_xor50;
  assign MulDiv_xor11 = MulDiv_xor23 ^ MulDiv_xor24;
  assign MulDiv_xor104 = mux_cond_60_pad ^ mux_cond_61_pad;
  assign MulDiv_xor51 = mux_cond_59_pad ^ MulDiv_xor104;
  assign MulDiv_xor106 = mux_cond_63_pad ^ mux_cond_64_pad;
  assign MulDiv_xor52 = mux_cond_62_pad ^ MulDiv_xor106;
  assign MulDiv_xor25 = MulDiv_xor51 ^ MulDiv_xor52;
  assign MulDiv_xor108 = mux_cond_66_pad ^ mux_cond_67_pad;
  assign MulDiv_xor53 = mux_cond_65_pad ^ MulDiv_xor108;
  assign MulDiv_xor109 = mux_cond_68_pad ^ mux_cond_69_pad;
  assign MulDiv_xor110 = mux_cond_70_pad ^ mux_cond_71_pad;
  assign MulDiv_xor54 = MulDiv_xor109 ^ MulDiv_xor110;
  assign MulDiv_xor26 = MulDiv_xor53 ^ MulDiv_xor54;
  assign MulDiv_xor12 = MulDiv_xor25 ^ MulDiv_xor26;
  assign MulDiv_xor5 = MulDiv_xor11 ^ MulDiv_xor12;
  assign MulDiv_xor112 = mux_cond_73_pad ^ mux_cond_74_pad;
  assign MulDiv_xor55 = mux_cond_72_pad ^ MulDiv_xor112;
  assign MulDiv_xor114 = mux_cond_76_pad ^ mux_cond_77_pad;
  assign MulDiv_xor56 = mux_cond_75_pad ^ MulDiv_xor114;
  assign MulDiv_xor27 = MulDiv_xor55 ^ MulDiv_xor56;
  assign MulDiv_xor116 = mux_cond_79_pad ^ mux_cond_80_pad;
  assign MulDiv_xor57 = mux_cond_78_pad ^ MulDiv_xor116;
  assign MulDiv_xor117 = mux_cond_81_pad ^ mux_cond_82_pad;
  assign MulDiv_xor118 = mux_cond_83_pad ^ mux_cond_84_pad;
  assign MulDiv_xor58 = MulDiv_xor117 ^ MulDiv_xor118;
  assign MulDiv_xor28 = MulDiv_xor57 ^ MulDiv_xor58;
  assign MulDiv_xor13 = MulDiv_xor27 ^ MulDiv_xor28;
  assign MulDiv_xor120 = mux_cond_86_pad ^ mux_cond_87_pad;
  assign MulDiv_xor59 = mux_cond_85_pad ^ MulDiv_xor120;
  assign MulDiv_xor122 = mux_cond_89_pad ^ mux_cond_90_pad;
  assign MulDiv_xor60 = mux_cond_88_pad ^ MulDiv_xor122;
  assign MulDiv_xor29 = MulDiv_xor59 ^ MulDiv_xor60;
  assign MulDiv_xor124 = mux_cond_92_pad ^ mux_cond_93_pad;
  assign MulDiv_xor61 = mux_cond_91_pad ^ MulDiv_xor124;
  assign MulDiv_xor125 = mux_cond_94_pad ^ mux_cond_95_pad;
  assign MulDiv_xor126 = mux_cond_96_pad ^ mux_cond_97_pad;
  assign MulDiv_xor62 = MulDiv_xor125 ^ MulDiv_xor126;
  assign MulDiv_xor30 = MulDiv_xor61 ^ MulDiv_xor62;
  assign MulDiv_xor14 = MulDiv_xor29 ^ MulDiv_xor30;
  assign MulDiv_xor6 = MulDiv_xor13 ^ MulDiv_xor14;
  assign MulDiv_xor2 = MulDiv_xor5 ^ MulDiv_xor6;
  assign MulDiv_xor0 = MulDiv_xor1 ^ MulDiv_xor2;
  assign io_covSum = MulDiv_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  req_dw = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  req_tag = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  count = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  neg_out = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  isHi = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  resHi = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {3{`RANDOM}};
  divisor = _RAND_7[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {5{`RANDOM}};
  remainder = _RAND_8[129:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  MulDiv_state = _RAND_9[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    MulDiv_cov[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  MulDiv_covSum = _RAND_11[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      state <= 3'h0;
    end else if (reset) begin
      state <= 3'h0;
    end else if (_T_448) begin
      if (cmdMul) begin
        state <= 3'h2;
      end else if (_T_449) begin
        state <= 3'h1;
      end else begin
        state <= 3'h3;
      end
    end else if (_T_447) begin
      state <= 3'h0;
    end else if (_T_100) begin
      if (_T_109) begin
        if (neg_out) begin
          state <= 3'h5;
        end else begin
          state <= 3'h7;
        end
      end else if (_T_48) begin
        if (_T_99) begin
          state <= 3'h6;
        end else if (_T_47) begin
          state <= 3'h7;
        end else if (_T_44) begin
          state <= 3'h3;
        end
      end else if (_T_47) begin
        state <= 3'h7;
      end else if (_T_44) begin
        state <= 3'h3;
      end
    end else if (_T_48) begin
      if (_T_99) begin
        state <= 3'h6;
      end else if (_T_47) begin
        state <= 3'h7;
      end else if (_T_44) begin
        state <= 3'h3;
      end
    end else if (_T_47) begin
      state <= 3'h7;
    end else if (_T_44) begin
      state <= 3'h3;
    end
    if (metaReset) begin
      req_dw <= 1'h0;
    end else if (_T_448) begin
      req_dw <= io_req_bits_dw;
    end
    if (metaReset) begin
      req_tag <= 5'h0;
    end else if (_T_448) begin
      req_tag <= io_req_bits_tag;
    end
    if (metaReset) begin
      count <= 7'h0;
    end else if (_T_448) begin
      count <= {{4'd0}, _T_455};
    end else if (_T_100) begin
      if (_T_440) begin
        count <= {{1'd0}, ~_T_434};
      end else begin
        count <= _T_97;
      end
    end else if (_T_48) begin
      count <= _T_97;
    end
    if (metaReset) begin
      neg_out <= 1'h0;
    end else if (_T_448) begin
      if (cmdHi) begin
        neg_out <= lhs_sign;
      end else begin
        neg_out <= _T_456;
      end
    end else if (_T_100) begin
      if (_T_445) begin
        neg_out <= 1'h0;
      end
    end
    if (metaReset) begin
      isHi <= 1'h0;
    end else if (_T_448) begin
      isHi <= cmdHi;
    end
    if (metaReset) begin
      resHi <= 1'h0;
    end else if (_T_448) begin
      resHi <= 1'h0;
    end else if (_T_100) begin
      if (_T_109) begin
        resHi <= isHi;
      end else if (_T_48) begin
        if (_T_99) begin
          resHi <= isHi;
        end else if (_T_47) begin
          resHi <= 1'h0;
        end
      end else if (_T_47) begin
        resHi <= 1'h0;
      end
    end else if (_T_48) begin
      if (_T_99) begin
        resHi <= isHi;
      end else if (_T_47) begin
        resHi <= 1'h0;
      end
    end else if (_T_47) begin
      resHi <= 1'h0;
    end
    if (metaReset) begin
      divisor <= 65'h0;
    end else if (_T_448) begin
      divisor <= _T_458;
    end else if (_T_44) begin
      if (divisor[63]) begin
        divisor <= subtractor;
      end
    end
    if (metaReset) begin
      remainder <= 130'h0;
    end else if (_T_448) begin
      remainder <= {{66'd0}, lhs_in};
    end else if (_T_100) begin
      remainder <= {{1'd0}, _GEN_16};
    end else if (_T_48) begin
      remainder <= _T_95;
    end else if (_T_47) begin
      remainder <= {{66'd0}, negated_remainder};
    end else if (_T_44) begin
      if (remainder[63]) begin
        remainder <= {{66'd0}, negated_remainder};
      end
    end
    MulDiv_state <= MulDiv_xor0;
    if (!(MulDiv_cov_read_data)) begin
      MulDiv_covSum <= MulDiv_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(MulDiv_cov_write_en & MulDiv_cov_write_mask) begin
      MulDiv_cov[MulDiv_cov_write_addr] <= MulDiv_cov_write_data; // @[Coverage map for MulDiv]
    end
  end
endmodule
module PlusArgTimeout(
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] PlusArgTimeout_covSum;
  assign PlusArgTimeout_covSum = 30'h0;
  assign io_covSum = PlusArgTimeout_covSum;
  assign metaAssert = 1'h0;
endmodule
module OptimizationBarrier(
  input  [19:0] io_x_ppn,
  input         io_x_u,
  input         io_x_ae,
  input         io_x_sw,
  input         io_x_sx,
  input         io_x_sr,
  input         io_x_pw,
  input         io_x_px,
  input         io_x_pr,
  input         io_x_ppp,
  input         io_x_pal,
  input         io_x_paa,
  input         io_x_eff,
  input         io_x_c,
  output [19:0] io_y_ppn,
  output        io_y_u,
  output        io_y_ae,
  output        io_y_sw,
  output        io_y_sx,
  output        io_y_sr,
  output        io_y_pw,
  output        io_y_px,
  output        io_y_pr,
  output        io_y_ppp,
  output        io_y_pal,
  output        io_y_paa,
  output        io_y_eff,
  output        io_y_c,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] OptimizationBarrier_covSum;
  assign io_y_ppn = io_x_ppn; // @[package.scala 241:12]
  assign io_y_u = io_x_u; // @[package.scala 241:12]
  assign io_y_ae = io_x_ae; // @[package.scala 241:12]
  assign io_y_sw = io_x_sw; // @[package.scala 241:12]
  assign io_y_sx = io_x_sx; // @[package.scala 241:12]
  assign io_y_sr = io_x_sr; // @[package.scala 241:12]
  assign io_y_pw = io_x_pw; // @[package.scala 241:12]
  assign io_y_px = io_x_px; // @[package.scala 241:12]
  assign io_y_pr = io_x_pr; // @[package.scala 241:12]
  assign io_y_ppp = io_x_ppp; // @[package.scala 241:12]
  assign io_y_pal = io_x_pal; // @[package.scala 241:12]
  assign io_y_paa = io_x_paa; // @[package.scala 241:12]
  assign io_y_eff = io_x_eff; // @[package.scala 241:12]
  assign io_y_c = io_x_c; // @[package.scala 241:12]
  assign OptimizationBarrier_covSum = 30'h0;
  assign io_covSum = OptimizationBarrier_covSum;
  assign metaAssert = 1'h0;
endmodule
module PMPChecker(
  input  [1:0]  io_prv,
  input         io_pmp_0_cfg_l,
  input  [1:0]  io_pmp_0_cfg_a,
  input         io_pmp_0_cfg_x,
  input         io_pmp_0_cfg_w,
  input         io_pmp_0_cfg_r,
  input  [29:0] io_pmp_0_addr,
  input  [31:0] io_pmp_0_mask,
  input         io_pmp_1_cfg_l,
  input  [1:0]  io_pmp_1_cfg_a,
  input         io_pmp_1_cfg_x,
  input         io_pmp_1_cfg_w,
  input         io_pmp_1_cfg_r,
  input  [29:0] io_pmp_1_addr,
  input  [31:0] io_pmp_1_mask,
  input         io_pmp_2_cfg_l,
  input  [1:0]  io_pmp_2_cfg_a,
  input         io_pmp_2_cfg_x,
  input         io_pmp_2_cfg_w,
  input         io_pmp_2_cfg_r,
  input  [29:0] io_pmp_2_addr,
  input  [31:0] io_pmp_2_mask,
  input         io_pmp_3_cfg_l,
  input  [1:0]  io_pmp_3_cfg_a,
  input         io_pmp_3_cfg_x,
  input         io_pmp_3_cfg_w,
  input         io_pmp_3_cfg_r,
  input  [29:0] io_pmp_3_addr,
  input  [31:0] io_pmp_3_mask,
  input         io_pmp_4_cfg_l,
  input  [1:0]  io_pmp_4_cfg_a,
  input         io_pmp_4_cfg_x,
  input         io_pmp_4_cfg_w,
  input         io_pmp_4_cfg_r,
  input  [29:0] io_pmp_4_addr,
  input  [31:0] io_pmp_4_mask,
  input         io_pmp_5_cfg_l,
  input  [1:0]  io_pmp_5_cfg_a,
  input         io_pmp_5_cfg_x,
  input         io_pmp_5_cfg_w,
  input         io_pmp_5_cfg_r,
  input  [29:0] io_pmp_5_addr,
  input  [31:0] io_pmp_5_mask,
  input         io_pmp_6_cfg_l,
  input  [1:0]  io_pmp_6_cfg_a,
  input         io_pmp_6_cfg_x,
  input         io_pmp_6_cfg_w,
  input         io_pmp_6_cfg_r,
  input  [29:0] io_pmp_6_addr,
  input  [31:0] io_pmp_6_mask,
  input         io_pmp_7_cfg_l,
  input  [1:0]  io_pmp_7_cfg_a,
  input         io_pmp_7_cfg_x,
  input         io_pmp_7_cfg_w,
  input         io_pmp_7_cfg_r,
  input  [29:0] io_pmp_7_addr,
  input  [31:0] io_pmp_7_mask,
  input  [31:0] io_addr,
  input  [1:0]  io_size,
  output        io_r,
  output        io_w,
  output        io_x,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  default_; // @[PMP.scala 157:56]
  wire [5:0] _T_3; // @[package.scala 212:77]
  wire [31:0] _GEN_0; // @[PMP.scala 70:26]
  wire [31:0] _T_6; // @[PMP.scala 70:26]
  wire [31:0] _T_8; // @[PMP.scala 62:36]
  wire [31:0] _T_10; // @[PMP.scala 62:48]
  wire [28:0] _T_12; // @[PMP.scala 71:53]
  wire [28:0] _T_14; // @[PMP.scala 65:47]
  wire [28:0] _T_16; // @[PMP.scala 65:52]
  wire  _T_17; // @[PMP.scala 65:58]
  wire [2:0] _T_23; // @[PMP.scala 72:55]
  wire [2:0] _T_25; // @[PMP.scala 65:47]
  wire [2:0] _T_27; // @[PMP.scala 65:52]
  wire  _T_28; // @[PMP.scala 65:58]
  wire  _T_29; // @[PMP.scala 73:16]
  wire [31:0] _T_36; // @[PMP.scala 62:36]
  wire [31:0] _T_38; // @[PMP.scala 62:48]
  wire [28:0] _T_40; // @[PMP.scala 82:52]
  wire  _T_41; // @[PMP.scala 82:39]
  wire [28:0] _T_48; // @[PMP.scala 83:41]
  wire  _T_49; // @[PMP.scala 83:69]
  wire [2:0] _T_51; // @[PMP.scala 84:42]
  wire [2:0] _T_56; // @[PMP.scala 84:64]
  wire  _T_57; // @[PMP.scala 84:53]
  wire  _T_58; // @[PMP.scala 85:30]
  wire  _T_59; // @[PMP.scala 85:16]
  wire  _T_67; // @[PMP.scala 82:39]
  wire  _T_75; // @[PMP.scala 83:69]
  wire  _T_83; // @[PMP.scala 84:53]
  wire  _T_84; // @[PMP.scala 85:30]
  wire  _T_85; // @[PMP.scala 85:16]
  wire  _T_86; // @[PMP.scala 96:48]
  wire  _T_87; // @[PMP.scala 134:61]
  wire  _T_88; // @[PMP.scala 134:8]
  wire  _T_90; // @[PMP.scala 165:26]
  wire [2:0] _T_110; // @[PMP.scala 125:123]
  wire  _T_111; // @[PMP.scala 125:145]
  wire  _T_112; // @[PMP.scala 125:88]
  wire [2:0] _T_128; // @[PMP.scala 126:113]
  wire  _T_129; // @[PMP.scala 126:146]
  wire  _T_130; // @[PMP.scala 126:83]
  wire  _T_131; // @[PMP.scala 127:46]
  wire [2:0] _T_135; // @[PMP.scala 128:32]
  wire  _T_136; // @[PMP.scala 128:57]
  wire  _T_138; // @[PMP.scala 129:8]
  wire  _T_190; // @[PMP.scala 183:40]
  wire  _T_191; // @[PMP.scala 183:26]
  wire  _T_192; // @[PMP.scala 184:40]
  wire  _T_193; // @[PMP.scala 184:26]
  wire  _T_194; // @[PMP.scala 185:40]
  wire  _T_195; // @[PMP.scala 185:26]
  wire  _T_196_cfg_x; // @[PMP.scala 186:8]
  wire  _T_196_cfg_w; // @[PMP.scala 186:8]
  wire  _T_196_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_202; // @[PMP.scala 70:26]
  wire [28:0] _T_212; // @[PMP.scala 65:52]
  wire  _T_213; // @[PMP.scala 65:58]
  wire [2:0] _T_221; // @[PMP.scala 65:47]
  wire [2:0] _T_223; // @[PMP.scala 65:52]
  wire  _T_224; // @[PMP.scala 65:58]
  wire  _T_225; // @[PMP.scala 73:16]
  wire [31:0] _T_232; // @[PMP.scala 62:36]
  wire [31:0] _T_234; // @[PMP.scala 62:48]
  wire [28:0] _T_236; // @[PMP.scala 82:52]
  wire  _T_237; // @[PMP.scala 82:39]
  wire [28:0] _T_244; // @[PMP.scala 83:41]
  wire  _T_245; // @[PMP.scala 83:69]
  wire [2:0] _T_252; // @[PMP.scala 84:64]
  wire  _T_253; // @[PMP.scala 84:53]
  wire  _T_254; // @[PMP.scala 85:30]
  wire  _T_255; // @[PMP.scala 85:16]
  wire  _T_279; // @[PMP.scala 84:53]
  wire  _T_280; // @[PMP.scala 85:30]
  wire  _T_281; // @[PMP.scala 85:16]
  wire  _T_282; // @[PMP.scala 96:48]
  wire  _T_283; // @[PMP.scala 134:61]
  wire  _T_284; // @[PMP.scala 134:8]
  wire  _T_286; // @[PMP.scala 165:26]
  wire [2:0] _T_306; // @[PMP.scala 125:123]
  wire  _T_307; // @[PMP.scala 125:145]
  wire  _T_308; // @[PMP.scala 125:88]
  wire [2:0] _T_324; // @[PMP.scala 126:113]
  wire  _T_325; // @[PMP.scala 126:146]
  wire  _T_326; // @[PMP.scala 126:83]
  wire  _T_327; // @[PMP.scala 127:46]
  wire [2:0] _T_331; // @[PMP.scala 128:32]
  wire  _T_332; // @[PMP.scala 128:57]
  wire  _T_334; // @[PMP.scala 129:8]
  wire  _T_386; // @[PMP.scala 183:40]
  wire  _T_387; // @[PMP.scala 183:26]
  wire  _T_388; // @[PMP.scala 184:40]
  wire  _T_389; // @[PMP.scala 184:26]
  wire  _T_390; // @[PMP.scala 185:40]
  wire  _T_391; // @[PMP.scala 185:26]
  wire  _T_392_cfg_x; // @[PMP.scala 186:8]
  wire  _T_392_cfg_w; // @[PMP.scala 186:8]
  wire  _T_392_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_398; // @[PMP.scala 70:26]
  wire [28:0] _T_408; // @[PMP.scala 65:52]
  wire  _T_409; // @[PMP.scala 65:58]
  wire [2:0] _T_417; // @[PMP.scala 65:47]
  wire [2:0] _T_419; // @[PMP.scala 65:52]
  wire  _T_420; // @[PMP.scala 65:58]
  wire  _T_421; // @[PMP.scala 73:16]
  wire [31:0] _T_428; // @[PMP.scala 62:36]
  wire [31:0] _T_430; // @[PMP.scala 62:48]
  wire [28:0] _T_432; // @[PMP.scala 82:52]
  wire  _T_433; // @[PMP.scala 82:39]
  wire [28:0] _T_440; // @[PMP.scala 83:41]
  wire  _T_441; // @[PMP.scala 83:69]
  wire [2:0] _T_448; // @[PMP.scala 84:64]
  wire  _T_449; // @[PMP.scala 84:53]
  wire  _T_450; // @[PMP.scala 85:30]
  wire  _T_451; // @[PMP.scala 85:16]
  wire  _T_475; // @[PMP.scala 84:53]
  wire  _T_476; // @[PMP.scala 85:30]
  wire  _T_477; // @[PMP.scala 85:16]
  wire  _T_478; // @[PMP.scala 96:48]
  wire  _T_479; // @[PMP.scala 134:61]
  wire  _T_480; // @[PMP.scala 134:8]
  wire  _T_482; // @[PMP.scala 165:26]
  wire [2:0] _T_502; // @[PMP.scala 125:123]
  wire  _T_503; // @[PMP.scala 125:145]
  wire  _T_504; // @[PMP.scala 125:88]
  wire [2:0] _T_520; // @[PMP.scala 126:113]
  wire  _T_521; // @[PMP.scala 126:146]
  wire  _T_522; // @[PMP.scala 126:83]
  wire  _T_523; // @[PMP.scala 127:46]
  wire [2:0] _T_527; // @[PMP.scala 128:32]
  wire  _T_528; // @[PMP.scala 128:57]
  wire  _T_530; // @[PMP.scala 129:8]
  wire  _T_582; // @[PMP.scala 183:40]
  wire  _T_583; // @[PMP.scala 183:26]
  wire  _T_584; // @[PMP.scala 184:40]
  wire  _T_585; // @[PMP.scala 184:26]
  wire  _T_586; // @[PMP.scala 185:40]
  wire  _T_587; // @[PMP.scala 185:26]
  wire  _T_588_cfg_x; // @[PMP.scala 186:8]
  wire  _T_588_cfg_w; // @[PMP.scala 186:8]
  wire  _T_588_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_594; // @[PMP.scala 70:26]
  wire [28:0] _T_604; // @[PMP.scala 65:52]
  wire  _T_605; // @[PMP.scala 65:58]
  wire [2:0] _T_613; // @[PMP.scala 65:47]
  wire [2:0] _T_615; // @[PMP.scala 65:52]
  wire  _T_616; // @[PMP.scala 65:58]
  wire  _T_617; // @[PMP.scala 73:16]
  wire [31:0] _T_624; // @[PMP.scala 62:36]
  wire [31:0] _T_626; // @[PMP.scala 62:48]
  wire [28:0] _T_628; // @[PMP.scala 82:52]
  wire  _T_629; // @[PMP.scala 82:39]
  wire [28:0] _T_636; // @[PMP.scala 83:41]
  wire  _T_637; // @[PMP.scala 83:69]
  wire [2:0] _T_644; // @[PMP.scala 84:64]
  wire  _T_645; // @[PMP.scala 84:53]
  wire  _T_646; // @[PMP.scala 85:30]
  wire  _T_647; // @[PMP.scala 85:16]
  wire  _T_671; // @[PMP.scala 84:53]
  wire  _T_672; // @[PMP.scala 85:30]
  wire  _T_673; // @[PMP.scala 85:16]
  wire  _T_674; // @[PMP.scala 96:48]
  wire  _T_675; // @[PMP.scala 134:61]
  wire  _T_676; // @[PMP.scala 134:8]
  wire  _T_678; // @[PMP.scala 165:26]
  wire [2:0] _T_698; // @[PMP.scala 125:123]
  wire  _T_699; // @[PMP.scala 125:145]
  wire  _T_700; // @[PMP.scala 125:88]
  wire [2:0] _T_716; // @[PMP.scala 126:113]
  wire  _T_717; // @[PMP.scala 126:146]
  wire  _T_718; // @[PMP.scala 126:83]
  wire  _T_719; // @[PMP.scala 127:46]
  wire [2:0] _T_723; // @[PMP.scala 128:32]
  wire  _T_724; // @[PMP.scala 128:57]
  wire  _T_726; // @[PMP.scala 129:8]
  wire  _T_778; // @[PMP.scala 183:40]
  wire  _T_779; // @[PMP.scala 183:26]
  wire  _T_780; // @[PMP.scala 184:40]
  wire  _T_781; // @[PMP.scala 184:26]
  wire  _T_782; // @[PMP.scala 185:40]
  wire  _T_783; // @[PMP.scala 185:26]
  wire  _T_784_cfg_x; // @[PMP.scala 186:8]
  wire  _T_784_cfg_w; // @[PMP.scala 186:8]
  wire  _T_784_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_790; // @[PMP.scala 70:26]
  wire [28:0] _T_800; // @[PMP.scala 65:52]
  wire  _T_801; // @[PMP.scala 65:58]
  wire [2:0] _T_809; // @[PMP.scala 65:47]
  wire [2:0] _T_811; // @[PMP.scala 65:52]
  wire  _T_812; // @[PMP.scala 65:58]
  wire  _T_813; // @[PMP.scala 73:16]
  wire [31:0] _T_820; // @[PMP.scala 62:36]
  wire [31:0] _T_822; // @[PMP.scala 62:48]
  wire [28:0] _T_824; // @[PMP.scala 82:52]
  wire  _T_825; // @[PMP.scala 82:39]
  wire [28:0] _T_832; // @[PMP.scala 83:41]
  wire  _T_833; // @[PMP.scala 83:69]
  wire [2:0] _T_840; // @[PMP.scala 84:64]
  wire  _T_841; // @[PMP.scala 84:53]
  wire  _T_842; // @[PMP.scala 85:30]
  wire  _T_843; // @[PMP.scala 85:16]
  wire  _T_867; // @[PMP.scala 84:53]
  wire  _T_868; // @[PMP.scala 85:30]
  wire  _T_869; // @[PMP.scala 85:16]
  wire  _T_870; // @[PMP.scala 96:48]
  wire  _T_871; // @[PMP.scala 134:61]
  wire  _T_872; // @[PMP.scala 134:8]
  wire  _T_874; // @[PMP.scala 165:26]
  wire [2:0] _T_894; // @[PMP.scala 125:123]
  wire  _T_895; // @[PMP.scala 125:145]
  wire  _T_896; // @[PMP.scala 125:88]
  wire [2:0] _T_912; // @[PMP.scala 126:113]
  wire  _T_913; // @[PMP.scala 126:146]
  wire  _T_914; // @[PMP.scala 126:83]
  wire  _T_915; // @[PMP.scala 127:46]
  wire [2:0] _T_919; // @[PMP.scala 128:32]
  wire  _T_920; // @[PMP.scala 128:57]
  wire  _T_922; // @[PMP.scala 129:8]
  wire  _T_974; // @[PMP.scala 183:40]
  wire  _T_975; // @[PMP.scala 183:26]
  wire  _T_976; // @[PMP.scala 184:40]
  wire  _T_977; // @[PMP.scala 184:26]
  wire  _T_978; // @[PMP.scala 185:40]
  wire  _T_979; // @[PMP.scala 185:26]
  wire  _T_980_cfg_x; // @[PMP.scala 186:8]
  wire  _T_980_cfg_w; // @[PMP.scala 186:8]
  wire  _T_980_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_986; // @[PMP.scala 70:26]
  wire [28:0] _T_996; // @[PMP.scala 65:52]
  wire  _T_997; // @[PMP.scala 65:58]
  wire [2:0] _T_1005; // @[PMP.scala 65:47]
  wire [2:0] _T_1007; // @[PMP.scala 65:52]
  wire  _T_1008; // @[PMP.scala 65:58]
  wire  _T_1009; // @[PMP.scala 73:16]
  wire [31:0] _T_1016; // @[PMP.scala 62:36]
  wire [31:0] _T_1018; // @[PMP.scala 62:48]
  wire [28:0] _T_1020; // @[PMP.scala 82:52]
  wire  _T_1021; // @[PMP.scala 82:39]
  wire [28:0] _T_1028; // @[PMP.scala 83:41]
  wire  _T_1029; // @[PMP.scala 83:69]
  wire [2:0] _T_1036; // @[PMP.scala 84:64]
  wire  _T_1037; // @[PMP.scala 84:53]
  wire  _T_1038; // @[PMP.scala 85:30]
  wire  _T_1039; // @[PMP.scala 85:16]
  wire  _T_1063; // @[PMP.scala 84:53]
  wire  _T_1064; // @[PMP.scala 85:30]
  wire  _T_1065; // @[PMP.scala 85:16]
  wire  _T_1066; // @[PMP.scala 96:48]
  wire  _T_1067; // @[PMP.scala 134:61]
  wire  _T_1068; // @[PMP.scala 134:8]
  wire  _T_1070; // @[PMP.scala 165:26]
  wire [2:0] _T_1090; // @[PMP.scala 125:123]
  wire  _T_1091; // @[PMP.scala 125:145]
  wire  _T_1092; // @[PMP.scala 125:88]
  wire [2:0] _T_1108; // @[PMP.scala 126:113]
  wire  _T_1109; // @[PMP.scala 126:146]
  wire  _T_1110; // @[PMP.scala 126:83]
  wire  _T_1111; // @[PMP.scala 127:46]
  wire [2:0] _T_1115; // @[PMP.scala 128:32]
  wire  _T_1116; // @[PMP.scala 128:57]
  wire  _T_1118; // @[PMP.scala 129:8]
  wire  _T_1170; // @[PMP.scala 183:40]
  wire  _T_1171; // @[PMP.scala 183:26]
  wire  _T_1172; // @[PMP.scala 184:40]
  wire  _T_1173; // @[PMP.scala 184:26]
  wire  _T_1174; // @[PMP.scala 185:40]
  wire  _T_1175; // @[PMP.scala 185:26]
  wire  _T_1176_cfg_x; // @[PMP.scala 186:8]
  wire  _T_1176_cfg_w; // @[PMP.scala 186:8]
  wire  _T_1176_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_1182; // @[PMP.scala 70:26]
  wire [28:0] _T_1192; // @[PMP.scala 65:52]
  wire  _T_1193; // @[PMP.scala 65:58]
  wire [2:0] _T_1201; // @[PMP.scala 65:47]
  wire [2:0] _T_1203; // @[PMP.scala 65:52]
  wire  _T_1204; // @[PMP.scala 65:58]
  wire  _T_1205; // @[PMP.scala 73:16]
  wire [31:0] _T_1212; // @[PMP.scala 62:36]
  wire [31:0] _T_1214; // @[PMP.scala 62:48]
  wire [28:0] _T_1216; // @[PMP.scala 82:52]
  wire  _T_1217; // @[PMP.scala 82:39]
  wire [28:0] _T_1224; // @[PMP.scala 83:41]
  wire  _T_1225; // @[PMP.scala 83:69]
  wire [2:0] _T_1232; // @[PMP.scala 84:64]
  wire  _T_1233; // @[PMP.scala 84:53]
  wire  _T_1234; // @[PMP.scala 85:30]
  wire  _T_1235; // @[PMP.scala 85:16]
  wire  _T_1259; // @[PMP.scala 84:53]
  wire  _T_1260; // @[PMP.scala 85:30]
  wire  _T_1261; // @[PMP.scala 85:16]
  wire  _T_1262; // @[PMP.scala 96:48]
  wire  _T_1263; // @[PMP.scala 134:61]
  wire  _T_1264; // @[PMP.scala 134:8]
  wire  _T_1266; // @[PMP.scala 165:26]
  wire [2:0] _T_1286; // @[PMP.scala 125:123]
  wire  _T_1287; // @[PMP.scala 125:145]
  wire  _T_1288; // @[PMP.scala 125:88]
  wire [2:0] _T_1304; // @[PMP.scala 126:113]
  wire  _T_1305; // @[PMP.scala 126:146]
  wire  _T_1306; // @[PMP.scala 126:83]
  wire  _T_1307; // @[PMP.scala 127:46]
  wire [2:0] _T_1311; // @[PMP.scala 128:32]
  wire  _T_1312; // @[PMP.scala 128:57]
  wire  _T_1314; // @[PMP.scala 129:8]
  wire  _T_1366; // @[PMP.scala 183:40]
  wire  _T_1367; // @[PMP.scala 183:26]
  wire  _T_1368; // @[PMP.scala 184:40]
  wire  _T_1369; // @[PMP.scala 184:26]
  wire  _T_1370; // @[PMP.scala 185:40]
  wire  _T_1371; // @[PMP.scala 185:26]
  wire  _T_1372_cfg_x; // @[PMP.scala 186:8]
  wire  _T_1372_cfg_w; // @[PMP.scala 186:8]
  wire  _T_1372_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_1378; // @[PMP.scala 70:26]
  wire [28:0] _T_1388; // @[PMP.scala 65:52]
  wire  _T_1389; // @[PMP.scala 65:58]
  wire [2:0] _T_1397; // @[PMP.scala 65:47]
  wire [2:0] _T_1399; // @[PMP.scala 65:52]
  wire  _T_1400; // @[PMP.scala 65:58]
  wire  _T_1401; // @[PMP.scala 73:16]
  wire  _T_1455; // @[PMP.scala 84:53]
  wire  _T_1456; // @[PMP.scala 85:30]
  wire  _T_1457; // @[PMP.scala 85:16]
  wire  _T_1459; // @[PMP.scala 134:61]
  wire  _T_1460; // @[PMP.scala 134:8]
  wire  _T_1462; // @[PMP.scala 165:26]
  wire [2:0] _T_1500; // @[PMP.scala 126:113]
  wire  _T_1501; // @[PMP.scala 126:146]
  wire  _T_1502; // @[PMP.scala 126:83]
  wire [2:0] _T_1507; // @[PMP.scala 128:32]
  wire  _T_1508; // @[PMP.scala 128:57]
  wire  _T_1510; // @[PMP.scala 129:8]
  wire  _T_1562; // @[PMP.scala 183:40]
  wire  _T_1563; // @[PMP.scala 183:26]
  wire  _T_1564; // @[PMP.scala 184:40]
  wire  _T_1565; // @[PMP.scala 184:26]
  wire  _T_1566; // @[PMP.scala 185:40]
  wire  _T_1567; // @[PMP.scala 185:26]
  wire [29:0] PMPChecker_covSum;
  assign default_ = io_prv > 2'h1; // @[PMP.scala 157:56]
  assign _T_3 = 6'h7 << io_size; // @[package.scala 212:77]
  assign _GEN_0 = {{29'd0}, ~_T_3[2:0]}; // @[PMP.scala 70:26]
  assign _T_6 = io_pmp_7_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _T_8 = {io_pmp_7_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_10 = ~_T_8 | 32'h3; // @[PMP.scala 62:48]
  assign _T_12 = ~_T_10[31:3]; // @[PMP.scala 71:53]
  assign _T_14 = io_addr[31:3] ^ _T_12; // @[PMP.scala 65:47]
  assign _T_16 = _T_14 & ~io_pmp_7_mask[31:3]; // @[PMP.scala 65:52]
  assign _T_17 = _T_16 == 29'h0; // @[PMP.scala 65:58]
  assign _T_23 = ~_T_10[2:0]; // @[PMP.scala 72:55]
  assign _T_25 = io_addr[2:0] ^ _T_23; // @[PMP.scala 65:47]
  assign _T_27 = _T_25 & ~_T_6[2:0]; // @[PMP.scala 65:52]
  assign _T_28 = _T_27 == 3'h0; // @[PMP.scala 65:58]
  assign _T_29 = _T_17 & _T_28; // @[PMP.scala 73:16]
  assign _T_36 = {io_pmp_6_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_38 = ~_T_36 | 32'h3; // @[PMP.scala 62:48]
  assign _T_40 = ~_T_38[31:3]; // @[PMP.scala 82:52]
  assign _T_41 = io_addr[31:3] < _T_40; // @[PMP.scala 82:39]
  assign _T_48 = io_addr[31:3] ^ _T_40; // @[PMP.scala 83:41]
  assign _T_49 = _T_48 == 29'h0; // @[PMP.scala 83:69]
  assign _T_51 = io_addr[2:0] | ~_T_3[2:0]; // @[PMP.scala 84:42]
  assign _T_56 = ~_T_38[2:0]; // @[PMP.scala 84:64]
  assign _T_57 = _T_51 < _T_56; // @[PMP.scala 84:53]
  assign _T_58 = _T_49 & _T_57; // @[PMP.scala 85:30]
  assign _T_59 = _T_41 | _T_58; // @[PMP.scala 85:16]
  assign _T_67 = io_addr[31:3] < _T_12; // @[PMP.scala 82:39]
  assign _T_75 = _T_14 == 29'h0; // @[PMP.scala 83:69]
  assign _T_83 = io_addr[2:0] < _T_23; // @[PMP.scala 84:53]
  assign _T_84 = _T_75 & _T_83; // @[PMP.scala 85:30]
  assign _T_85 = _T_67 | _T_84; // @[PMP.scala 85:16]
  assign _T_86 = ~_T_59 & _T_85; // @[PMP.scala 96:48]
  assign _T_87 = io_pmp_7_cfg_a[0] & _T_86; // @[PMP.scala 134:61]
  assign _T_88 = io_pmp_7_cfg_a[1] ? _T_29 : _T_87; // @[PMP.scala 134:8]
  assign _T_90 = default_ & ~io_pmp_7_cfg_l; // @[PMP.scala 165:26]
  assign _T_110 = _T_56 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _T_111 = _T_110 != 3'h0; // @[PMP.scala 125:145]
  assign _T_112 = _T_49 & _T_111; // @[PMP.scala 125:88]
  assign _T_128 = _T_23 & _T_51; // @[PMP.scala 126:113]
  assign _T_129 = _T_128 != 3'h0; // @[PMP.scala 126:146]
  assign _T_130 = _T_75 & _T_129; // @[PMP.scala 126:83]
  assign _T_131 = _T_112 | _T_130; // @[PMP.scala 127:46]
  assign _T_135 = ~_T_3[2:0] & ~io_pmp_7_mask[2:0]; // @[PMP.scala 128:32]
  assign _T_136 = _T_135 == 3'h0; // @[PMP.scala 128:57]
  assign _T_138 = io_pmp_7_cfg_a[1] ? _T_136 : ~_T_131; // @[PMP.scala 129:8]
  assign _T_190 = io_pmp_7_cfg_r | _T_90; // @[PMP.scala 183:40]
  assign _T_191 = _T_138 & _T_190; // @[PMP.scala 183:26]
  assign _T_192 = io_pmp_7_cfg_w | _T_90; // @[PMP.scala 184:40]
  assign _T_193 = _T_138 & _T_192; // @[PMP.scala 184:26]
  assign _T_194 = io_pmp_7_cfg_x | _T_90; // @[PMP.scala 185:40]
  assign _T_195 = _T_138 & _T_194; // @[PMP.scala 185:26]
  assign _T_196_cfg_x = _T_88 ? _T_195 : default_; // @[PMP.scala 186:8]
  assign _T_196_cfg_w = _T_88 ? _T_193 : default_; // @[PMP.scala 186:8]
  assign _T_196_cfg_r = _T_88 ? _T_191 : default_; // @[PMP.scala 186:8]
  assign _T_202 = io_pmp_6_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _T_212 = _T_48 & ~io_pmp_6_mask[31:3]; // @[PMP.scala 65:52]
  assign _T_213 = _T_212 == 29'h0; // @[PMP.scala 65:58]
  assign _T_221 = io_addr[2:0] ^ _T_56; // @[PMP.scala 65:47]
  assign _T_223 = _T_221 & ~_T_202[2:0]; // @[PMP.scala 65:52]
  assign _T_224 = _T_223 == 3'h0; // @[PMP.scala 65:58]
  assign _T_225 = _T_213 & _T_224; // @[PMP.scala 73:16]
  assign _T_232 = {io_pmp_5_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_234 = ~_T_232 | 32'h3; // @[PMP.scala 62:48]
  assign _T_236 = ~_T_234[31:3]; // @[PMP.scala 82:52]
  assign _T_237 = io_addr[31:3] < _T_236; // @[PMP.scala 82:39]
  assign _T_244 = io_addr[31:3] ^ _T_236; // @[PMP.scala 83:41]
  assign _T_245 = _T_244 == 29'h0; // @[PMP.scala 83:69]
  assign _T_252 = ~_T_234[2:0]; // @[PMP.scala 84:64]
  assign _T_253 = _T_51 < _T_252; // @[PMP.scala 84:53]
  assign _T_254 = _T_245 & _T_253; // @[PMP.scala 85:30]
  assign _T_255 = _T_237 | _T_254; // @[PMP.scala 85:16]
  assign _T_279 = io_addr[2:0] < _T_56; // @[PMP.scala 84:53]
  assign _T_280 = _T_49 & _T_279; // @[PMP.scala 85:30]
  assign _T_281 = _T_41 | _T_280; // @[PMP.scala 85:16]
  assign _T_282 = ~_T_255 & _T_281; // @[PMP.scala 96:48]
  assign _T_283 = io_pmp_6_cfg_a[0] & _T_282; // @[PMP.scala 134:61]
  assign _T_284 = io_pmp_6_cfg_a[1] ? _T_225 : _T_283; // @[PMP.scala 134:8]
  assign _T_286 = default_ & ~io_pmp_6_cfg_l; // @[PMP.scala 165:26]
  assign _T_306 = _T_252 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _T_307 = _T_306 != 3'h0; // @[PMP.scala 125:145]
  assign _T_308 = _T_245 & _T_307; // @[PMP.scala 125:88]
  assign _T_324 = _T_56 & _T_51; // @[PMP.scala 126:113]
  assign _T_325 = _T_324 != 3'h0; // @[PMP.scala 126:146]
  assign _T_326 = _T_49 & _T_325; // @[PMP.scala 126:83]
  assign _T_327 = _T_308 | _T_326; // @[PMP.scala 127:46]
  assign _T_331 = ~_T_3[2:0] & ~io_pmp_6_mask[2:0]; // @[PMP.scala 128:32]
  assign _T_332 = _T_331 == 3'h0; // @[PMP.scala 128:57]
  assign _T_334 = io_pmp_6_cfg_a[1] ? _T_332 : ~_T_327; // @[PMP.scala 129:8]
  assign _T_386 = io_pmp_6_cfg_r | _T_286; // @[PMP.scala 183:40]
  assign _T_387 = _T_334 & _T_386; // @[PMP.scala 183:26]
  assign _T_388 = io_pmp_6_cfg_w | _T_286; // @[PMP.scala 184:40]
  assign _T_389 = _T_334 & _T_388; // @[PMP.scala 184:26]
  assign _T_390 = io_pmp_6_cfg_x | _T_286; // @[PMP.scala 185:40]
  assign _T_391 = _T_334 & _T_390; // @[PMP.scala 185:26]
  assign _T_392_cfg_x = _T_284 ? _T_391 : _T_196_cfg_x; // @[PMP.scala 186:8]
  assign _T_392_cfg_w = _T_284 ? _T_389 : _T_196_cfg_w; // @[PMP.scala 186:8]
  assign _T_392_cfg_r = _T_284 ? _T_387 : _T_196_cfg_r; // @[PMP.scala 186:8]
  assign _T_398 = io_pmp_5_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _T_408 = _T_244 & ~io_pmp_5_mask[31:3]; // @[PMP.scala 65:52]
  assign _T_409 = _T_408 == 29'h0; // @[PMP.scala 65:58]
  assign _T_417 = io_addr[2:0] ^ _T_252; // @[PMP.scala 65:47]
  assign _T_419 = _T_417 & ~_T_398[2:0]; // @[PMP.scala 65:52]
  assign _T_420 = _T_419 == 3'h0; // @[PMP.scala 65:58]
  assign _T_421 = _T_409 & _T_420; // @[PMP.scala 73:16]
  assign _T_428 = {io_pmp_4_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_430 = ~_T_428 | 32'h3; // @[PMP.scala 62:48]
  assign _T_432 = ~_T_430[31:3]; // @[PMP.scala 82:52]
  assign _T_433 = io_addr[31:3] < _T_432; // @[PMP.scala 82:39]
  assign _T_440 = io_addr[31:3] ^ _T_432; // @[PMP.scala 83:41]
  assign _T_441 = _T_440 == 29'h0; // @[PMP.scala 83:69]
  assign _T_448 = ~_T_430[2:0]; // @[PMP.scala 84:64]
  assign _T_449 = _T_51 < _T_448; // @[PMP.scala 84:53]
  assign _T_450 = _T_441 & _T_449; // @[PMP.scala 85:30]
  assign _T_451 = _T_433 | _T_450; // @[PMP.scala 85:16]
  assign _T_475 = io_addr[2:0] < _T_252; // @[PMP.scala 84:53]
  assign _T_476 = _T_245 & _T_475; // @[PMP.scala 85:30]
  assign _T_477 = _T_237 | _T_476; // @[PMP.scala 85:16]
  assign _T_478 = ~_T_451 & _T_477; // @[PMP.scala 96:48]
  assign _T_479 = io_pmp_5_cfg_a[0] & _T_478; // @[PMP.scala 134:61]
  assign _T_480 = io_pmp_5_cfg_a[1] ? _T_421 : _T_479; // @[PMP.scala 134:8]
  assign _T_482 = default_ & ~io_pmp_5_cfg_l; // @[PMP.scala 165:26]
  assign _T_502 = _T_448 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _T_503 = _T_502 != 3'h0; // @[PMP.scala 125:145]
  assign _T_504 = _T_441 & _T_503; // @[PMP.scala 125:88]
  assign _T_520 = _T_252 & _T_51; // @[PMP.scala 126:113]
  assign _T_521 = _T_520 != 3'h0; // @[PMP.scala 126:146]
  assign _T_522 = _T_245 & _T_521; // @[PMP.scala 126:83]
  assign _T_523 = _T_504 | _T_522; // @[PMP.scala 127:46]
  assign _T_527 = ~_T_3[2:0] & ~io_pmp_5_mask[2:0]; // @[PMP.scala 128:32]
  assign _T_528 = _T_527 == 3'h0; // @[PMP.scala 128:57]
  assign _T_530 = io_pmp_5_cfg_a[1] ? _T_528 : ~_T_523; // @[PMP.scala 129:8]
  assign _T_582 = io_pmp_5_cfg_r | _T_482; // @[PMP.scala 183:40]
  assign _T_583 = _T_530 & _T_582; // @[PMP.scala 183:26]
  assign _T_584 = io_pmp_5_cfg_w | _T_482; // @[PMP.scala 184:40]
  assign _T_585 = _T_530 & _T_584; // @[PMP.scala 184:26]
  assign _T_586 = io_pmp_5_cfg_x | _T_482; // @[PMP.scala 185:40]
  assign _T_587 = _T_530 & _T_586; // @[PMP.scala 185:26]
  assign _T_588_cfg_x = _T_480 ? _T_587 : _T_392_cfg_x; // @[PMP.scala 186:8]
  assign _T_588_cfg_w = _T_480 ? _T_585 : _T_392_cfg_w; // @[PMP.scala 186:8]
  assign _T_588_cfg_r = _T_480 ? _T_583 : _T_392_cfg_r; // @[PMP.scala 186:8]
  assign _T_594 = io_pmp_4_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _T_604 = _T_440 & ~io_pmp_4_mask[31:3]; // @[PMP.scala 65:52]
  assign _T_605 = _T_604 == 29'h0; // @[PMP.scala 65:58]
  assign _T_613 = io_addr[2:0] ^ _T_448; // @[PMP.scala 65:47]
  assign _T_615 = _T_613 & ~_T_594[2:0]; // @[PMP.scala 65:52]
  assign _T_616 = _T_615 == 3'h0; // @[PMP.scala 65:58]
  assign _T_617 = _T_605 & _T_616; // @[PMP.scala 73:16]
  assign _T_624 = {io_pmp_3_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_626 = ~_T_624 | 32'h3; // @[PMP.scala 62:48]
  assign _T_628 = ~_T_626[31:3]; // @[PMP.scala 82:52]
  assign _T_629 = io_addr[31:3] < _T_628; // @[PMP.scala 82:39]
  assign _T_636 = io_addr[31:3] ^ _T_628; // @[PMP.scala 83:41]
  assign _T_637 = _T_636 == 29'h0; // @[PMP.scala 83:69]
  assign _T_644 = ~_T_626[2:0]; // @[PMP.scala 84:64]
  assign _T_645 = _T_51 < _T_644; // @[PMP.scala 84:53]
  assign _T_646 = _T_637 & _T_645; // @[PMP.scala 85:30]
  assign _T_647 = _T_629 | _T_646; // @[PMP.scala 85:16]
  assign _T_671 = io_addr[2:0] < _T_448; // @[PMP.scala 84:53]
  assign _T_672 = _T_441 & _T_671; // @[PMP.scala 85:30]
  assign _T_673 = _T_433 | _T_672; // @[PMP.scala 85:16]
  assign _T_674 = ~_T_647 & _T_673; // @[PMP.scala 96:48]
  assign _T_675 = io_pmp_4_cfg_a[0] & _T_674; // @[PMP.scala 134:61]
  assign _T_676 = io_pmp_4_cfg_a[1] ? _T_617 : _T_675; // @[PMP.scala 134:8]
  assign _T_678 = default_ & ~io_pmp_4_cfg_l; // @[PMP.scala 165:26]
  assign _T_698 = _T_644 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _T_699 = _T_698 != 3'h0; // @[PMP.scala 125:145]
  assign _T_700 = _T_637 & _T_699; // @[PMP.scala 125:88]
  assign _T_716 = _T_448 & _T_51; // @[PMP.scala 126:113]
  assign _T_717 = _T_716 != 3'h0; // @[PMP.scala 126:146]
  assign _T_718 = _T_441 & _T_717; // @[PMP.scala 126:83]
  assign _T_719 = _T_700 | _T_718; // @[PMP.scala 127:46]
  assign _T_723 = ~_T_3[2:0] & ~io_pmp_4_mask[2:0]; // @[PMP.scala 128:32]
  assign _T_724 = _T_723 == 3'h0; // @[PMP.scala 128:57]
  assign _T_726 = io_pmp_4_cfg_a[1] ? _T_724 : ~_T_719; // @[PMP.scala 129:8]
  assign _T_778 = io_pmp_4_cfg_r | _T_678; // @[PMP.scala 183:40]
  assign _T_779 = _T_726 & _T_778; // @[PMP.scala 183:26]
  assign _T_780 = io_pmp_4_cfg_w | _T_678; // @[PMP.scala 184:40]
  assign _T_781 = _T_726 & _T_780; // @[PMP.scala 184:26]
  assign _T_782 = io_pmp_4_cfg_x | _T_678; // @[PMP.scala 185:40]
  assign _T_783 = _T_726 & _T_782; // @[PMP.scala 185:26]
  assign _T_784_cfg_x = _T_676 ? _T_783 : _T_588_cfg_x; // @[PMP.scala 186:8]
  assign _T_784_cfg_w = _T_676 ? _T_781 : _T_588_cfg_w; // @[PMP.scala 186:8]
  assign _T_784_cfg_r = _T_676 ? _T_779 : _T_588_cfg_r; // @[PMP.scala 186:8]
  assign _T_790 = io_pmp_3_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _T_800 = _T_636 & ~io_pmp_3_mask[31:3]; // @[PMP.scala 65:52]
  assign _T_801 = _T_800 == 29'h0; // @[PMP.scala 65:58]
  assign _T_809 = io_addr[2:0] ^ _T_644; // @[PMP.scala 65:47]
  assign _T_811 = _T_809 & ~_T_790[2:0]; // @[PMP.scala 65:52]
  assign _T_812 = _T_811 == 3'h0; // @[PMP.scala 65:58]
  assign _T_813 = _T_801 & _T_812; // @[PMP.scala 73:16]
  assign _T_820 = {io_pmp_2_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_822 = ~_T_820 | 32'h3; // @[PMP.scala 62:48]
  assign _T_824 = ~_T_822[31:3]; // @[PMP.scala 82:52]
  assign _T_825 = io_addr[31:3] < _T_824; // @[PMP.scala 82:39]
  assign _T_832 = io_addr[31:3] ^ _T_824; // @[PMP.scala 83:41]
  assign _T_833 = _T_832 == 29'h0; // @[PMP.scala 83:69]
  assign _T_840 = ~_T_822[2:0]; // @[PMP.scala 84:64]
  assign _T_841 = _T_51 < _T_840; // @[PMP.scala 84:53]
  assign _T_842 = _T_833 & _T_841; // @[PMP.scala 85:30]
  assign _T_843 = _T_825 | _T_842; // @[PMP.scala 85:16]
  assign _T_867 = io_addr[2:0] < _T_644; // @[PMP.scala 84:53]
  assign _T_868 = _T_637 & _T_867; // @[PMP.scala 85:30]
  assign _T_869 = _T_629 | _T_868; // @[PMP.scala 85:16]
  assign _T_870 = ~_T_843 & _T_869; // @[PMP.scala 96:48]
  assign _T_871 = io_pmp_3_cfg_a[0] & _T_870; // @[PMP.scala 134:61]
  assign _T_872 = io_pmp_3_cfg_a[1] ? _T_813 : _T_871; // @[PMP.scala 134:8]
  assign _T_874 = default_ & ~io_pmp_3_cfg_l; // @[PMP.scala 165:26]
  assign _T_894 = _T_840 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _T_895 = _T_894 != 3'h0; // @[PMP.scala 125:145]
  assign _T_896 = _T_833 & _T_895; // @[PMP.scala 125:88]
  assign _T_912 = _T_644 & _T_51; // @[PMP.scala 126:113]
  assign _T_913 = _T_912 != 3'h0; // @[PMP.scala 126:146]
  assign _T_914 = _T_637 & _T_913; // @[PMP.scala 126:83]
  assign _T_915 = _T_896 | _T_914; // @[PMP.scala 127:46]
  assign _T_919 = ~_T_3[2:0] & ~io_pmp_3_mask[2:0]; // @[PMP.scala 128:32]
  assign _T_920 = _T_919 == 3'h0; // @[PMP.scala 128:57]
  assign _T_922 = io_pmp_3_cfg_a[1] ? _T_920 : ~_T_915; // @[PMP.scala 129:8]
  assign _T_974 = io_pmp_3_cfg_r | _T_874; // @[PMP.scala 183:40]
  assign _T_975 = _T_922 & _T_974; // @[PMP.scala 183:26]
  assign _T_976 = io_pmp_3_cfg_w | _T_874; // @[PMP.scala 184:40]
  assign _T_977 = _T_922 & _T_976; // @[PMP.scala 184:26]
  assign _T_978 = io_pmp_3_cfg_x | _T_874; // @[PMP.scala 185:40]
  assign _T_979 = _T_922 & _T_978; // @[PMP.scala 185:26]
  assign _T_980_cfg_x = _T_872 ? _T_979 : _T_784_cfg_x; // @[PMP.scala 186:8]
  assign _T_980_cfg_w = _T_872 ? _T_977 : _T_784_cfg_w; // @[PMP.scala 186:8]
  assign _T_980_cfg_r = _T_872 ? _T_975 : _T_784_cfg_r; // @[PMP.scala 186:8]
  assign _T_986 = io_pmp_2_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _T_996 = _T_832 & ~io_pmp_2_mask[31:3]; // @[PMP.scala 65:52]
  assign _T_997 = _T_996 == 29'h0; // @[PMP.scala 65:58]
  assign _T_1005 = io_addr[2:0] ^ _T_840; // @[PMP.scala 65:47]
  assign _T_1007 = _T_1005 & ~_T_986[2:0]; // @[PMP.scala 65:52]
  assign _T_1008 = _T_1007 == 3'h0; // @[PMP.scala 65:58]
  assign _T_1009 = _T_997 & _T_1008; // @[PMP.scala 73:16]
  assign _T_1016 = {io_pmp_1_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_1018 = ~_T_1016 | 32'h3; // @[PMP.scala 62:48]
  assign _T_1020 = ~_T_1018[31:3]; // @[PMP.scala 82:52]
  assign _T_1021 = io_addr[31:3] < _T_1020; // @[PMP.scala 82:39]
  assign _T_1028 = io_addr[31:3] ^ _T_1020; // @[PMP.scala 83:41]
  assign _T_1029 = _T_1028 == 29'h0; // @[PMP.scala 83:69]
  assign _T_1036 = ~_T_1018[2:0]; // @[PMP.scala 84:64]
  assign _T_1037 = _T_51 < _T_1036; // @[PMP.scala 84:53]
  assign _T_1038 = _T_1029 & _T_1037; // @[PMP.scala 85:30]
  assign _T_1039 = _T_1021 | _T_1038; // @[PMP.scala 85:16]
  assign _T_1063 = io_addr[2:0] < _T_840; // @[PMP.scala 84:53]
  assign _T_1064 = _T_833 & _T_1063; // @[PMP.scala 85:30]
  assign _T_1065 = _T_825 | _T_1064; // @[PMP.scala 85:16]
  assign _T_1066 = ~_T_1039 & _T_1065; // @[PMP.scala 96:48]
  assign _T_1067 = io_pmp_2_cfg_a[0] & _T_1066; // @[PMP.scala 134:61]
  assign _T_1068 = io_pmp_2_cfg_a[1] ? _T_1009 : _T_1067; // @[PMP.scala 134:8]
  assign _T_1070 = default_ & ~io_pmp_2_cfg_l; // @[PMP.scala 165:26]
  assign _T_1090 = _T_1036 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _T_1091 = _T_1090 != 3'h0; // @[PMP.scala 125:145]
  assign _T_1092 = _T_1029 & _T_1091; // @[PMP.scala 125:88]
  assign _T_1108 = _T_840 & _T_51; // @[PMP.scala 126:113]
  assign _T_1109 = _T_1108 != 3'h0; // @[PMP.scala 126:146]
  assign _T_1110 = _T_833 & _T_1109; // @[PMP.scala 126:83]
  assign _T_1111 = _T_1092 | _T_1110; // @[PMP.scala 127:46]
  assign _T_1115 = ~_T_3[2:0] & ~io_pmp_2_mask[2:0]; // @[PMP.scala 128:32]
  assign _T_1116 = _T_1115 == 3'h0; // @[PMP.scala 128:57]
  assign _T_1118 = io_pmp_2_cfg_a[1] ? _T_1116 : ~_T_1111; // @[PMP.scala 129:8]
  assign _T_1170 = io_pmp_2_cfg_r | _T_1070; // @[PMP.scala 183:40]
  assign _T_1171 = _T_1118 & _T_1170; // @[PMP.scala 183:26]
  assign _T_1172 = io_pmp_2_cfg_w | _T_1070; // @[PMP.scala 184:40]
  assign _T_1173 = _T_1118 & _T_1172; // @[PMP.scala 184:26]
  assign _T_1174 = io_pmp_2_cfg_x | _T_1070; // @[PMP.scala 185:40]
  assign _T_1175 = _T_1118 & _T_1174; // @[PMP.scala 185:26]
  assign _T_1176_cfg_x = _T_1068 ? _T_1175 : _T_980_cfg_x; // @[PMP.scala 186:8]
  assign _T_1176_cfg_w = _T_1068 ? _T_1173 : _T_980_cfg_w; // @[PMP.scala 186:8]
  assign _T_1176_cfg_r = _T_1068 ? _T_1171 : _T_980_cfg_r; // @[PMP.scala 186:8]
  assign _T_1182 = io_pmp_1_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _T_1192 = _T_1028 & ~io_pmp_1_mask[31:3]; // @[PMP.scala 65:52]
  assign _T_1193 = _T_1192 == 29'h0; // @[PMP.scala 65:58]
  assign _T_1201 = io_addr[2:0] ^ _T_1036; // @[PMP.scala 65:47]
  assign _T_1203 = _T_1201 & ~_T_1182[2:0]; // @[PMP.scala 65:52]
  assign _T_1204 = _T_1203 == 3'h0; // @[PMP.scala 65:58]
  assign _T_1205 = _T_1193 & _T_1204; // @[PMP.scala 73:16]
  assign _T_1212 = {io_pmp_0_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_1214 = ~_T_1212 | 32'h3; // @[PMP.scala 62:48]
  assign _T_1216 = ~_T_1214[31:3]; // @[PMP.scala 82:52]
  assign _T_1217 = io_addr[31:3] < _T_1216; // @[PMP.scala 82:39]
  assign _T_1224 = io_addr[31:3] ^ _T_1216; // @[PMP.scala 83:41]
  assign _T_1225 = _T_1224 == 29'h0; // @[PMP.scala 83:69]
  assign _T_1232 = ~_T_1214[2:0]; // @[PMP.scala 84:64]
  assign _T_1233 = _T_51 < _T_1232; // @[PMP.scala 84:53]
  assign _T_1234 = _T_1225 & _T_1233; // @[PMP.scala 85:30]
  assign _T_1235 = _T_1217 | _T_1234; // @[PMP.scala 85:16]
  assign _T_1259 = io_addr[2:0] < _T_1036; // @[PMP.scala 84:53]
  assign _T_1260 = _T_1029 & _T_1259; // @[PMP.scala 85:30]
  assign _T_1261 = _T_1021 | _T_1260; // @[PMP.scala 85:16]
  assign _T_1262 = ~_T_1235 & _T_1261; // @[PMP.scala 96:48]
  assign _T_1263 = io_pmp_1_cfg_a[0] & _T_1262; // @[PMP.scala 134:61]
  assign _T_1264 = io_pmp_1_cfg_a[1] ? _T_1205 : _T_1263; // @[PMP.scala 134:8]
  assign _T_1266 = default_ & ~io_pmp_1_cfg_l; // @[PMP.scala 165:26]
  assign _T_1286 = _T_1232 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _T_1287 = _T_1286 != 3'h0; // @[PMP.scala 125:145]
  assign _T_1288 = _T_1225 & _T_1287; // @[PMP.scala 125:88]
  assign _T_1304 = _T_1036 & _T_51; // @[PMP.scala 126:113]
  assign _T_1305 = _T_1304 != 3'h0; // @[PMP.scala 126:146]
  assign _T_1306 = _T_1029 & _T_1305; // @[PMP.scala 126:83]
  assign _T_1307 = _T_1288 | _T_1306; // @[PMP.scala 127:46]
  assign _T_1311 = ~_T_3[2:0] & ~io_pmp_1_mask[2:0]; // @[PMP.scala 128:32]
  assign _T_1312 = _T_1311 == 3'h0; // @[PMP.scala 128:57]
  assign _T_1314 = io_pmp_1_cfg_a[1] ? _T_1312 : ~_T_1307; // @[PMP.scala 129:8]
  assign _T_1366 = io_pmp_1_cfg_r | _T_1266; // @[PMP.scala 183:40]
  assign _T_1367 = _T_1314 & _T_1366; // @[PMP.scala 183:26]
  assign _T_1368 = io_pmp_1_cfg_w | _T_1266; // @[PMP.scala 184:40]
  assign _T_1369 = _T_1314 & _T_1368; // @[PMP.scala 184:26]
  assign _T_1370 = io_pmp_1_cfg_x | _T_1266; // @[PMP.scala 185:40]
  assign _T_1371 = _T_1314 & _T_1370; // @[PMP.scala 185:26]
  assign _T_1372_cfg_x = _T_1264 ? _T_1371 : _T_1176_cfg_x; // @[PMP.scala 186:8]
  assign _T_1372_cfg_w = _T_1264 ? _T_1369 : _T_1176_cfg_w; // @[PMP.scala 186:8]
  assign _T_1372_cfg_r = _T_1264 ? _T_1367 : _T_1176_cfg_r; // @[PMP.scala 186:8]
  assign _T_1378 = io_pmp_0_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _T_1388 = _T_1224 & ~io_pmp_0_mask[31:3]; // @[PMP.scala 65:52]
  assign _T_1389 = _T_1388 == 29'h0; // @[PMP.scala 65:58]
  assign _T_1397 = io_addr[2:0] ^ _T_1232; // @[PMP.scala 65:47]
  assign _T_1399 = _T_1397 & ~_T_1378[2:0]; // @[PMP.scala 65:52]
  assign _T_1400 = _T_1399 == 3'h0; // @[PMP.scala 65:58]
  assign _T_1401 = _T_1389 & _T_1400; // @[PMP.scala 73:16]
  assign _T_1455 = io_addr[2:0] < _T_1232; // @[PMP.scala 84:53]
  assign _T_1456 = _T_1225 & _T_1455; // @[PMP.scala 85:30]
  assign _T_1457 = _T_1217 | _T_1456; // @[PMP.scala 85:16]
  assign _T_1459 = io_pmp_0_cfg_a[0] & _T_1457; // @[PMP.scala 134:61]
  assign _T_1460 = io_pmp_0_cfg_a[1] ? _T_1401 : _T_1459; // @[PMP.scala 134:8]
  assign _T_1462 = default_ & ~io_pmp_0_cfg_l; // @[PMP.scala 165:26]
  assign _T_1500 = _T_1232 & _T_51; // @[PMP.scala 126:113]
  assign _T_1501 = _T_1500 != 3'h0; // @[PMP.scala 126:146]
  assign _T_1502 = _T_1225 & _T_1501; // @[PMP.scala 126:83]
  assign _T_1507 = ~_T_3[2:0] & ~io_pmp_0_mask[2:0]; // @[PMP.scala 128:32]
  assign _T_1508 = _T_1507 == 3'h0; // @[PMP.scala 128:57]
  assign _T_1510 = io_pmp_0_cfg_a[1] ? _T_1508 : ~_T_1502; // @[PMP.scala 129:8]
  assign _T_1562 = io_pmp_0_cfg_r | _T_1462; // @[PMP.scala 183:40]
  assign _T_1563 = _T_1510 & _T_1562; // @[PMP.scala 183:26]
  assign _T_1564 = io_pmp_0_cfg_w | _T_1462; // @[PMP.scala 184:40]
  assign _T_1565 = _T_1510 & _T_1564; // @[PMP.scala 184:26]
  assign _T_1566 = io_pmp_0_cfg_x | _T_1462; // @[PMP.scala 185:40]
  assign _T_1567 = _T_1510 & _T_1566; // @[PMP.scala 185:26]
  assign io_r = _T_1460 ? _T_1563 : _T_1372_cfg_r; // @[PMP.scala 189:8]
  assign io_w = _T_1460 ? _T_1565 : _T_1372_cfg_w; // @[PMP.scala 190:8]
  assign io_x = _T_1460 ? _T_1567 : _T_1372_cfg_x; // @[PMP.scala 191:8]
  assign PMPChecker_covSum = 30'h0;
  assign io_covSum = PMPChecker_covSum;
  assign metaAssert = 1'h0;
endmodule
module PMPChecker_2(
  input  [1:0]  io_prv,
  input         io_pmp_0_cfg_l,
  input  [1:0]  io_pmp_0_cfg_a,
  input         io_pmp_0_cfg_x,
  input         io_pmp_0_cfg_w,
  input         io_pmp_0_cfg_r,
  input  [29:0] io_pmp_0_addr,
  input  [31:0] io_pmp_0_mask,
  input         io_pmp_1_cfg_l,
  input  [1:0]  io_pmp_1_cfg_a,
  input         io_pmp_1_cfg_x,
  input         io_pmp_1_cfg_w,
  input         io_pmp_1_cfg_r,
  input  [29:0] io_pmp_1_addr,
  input  [31:0] io_pmp_1_mask,
  input         io_pmp_2_cfg_l,
  input  [1:0]  io_pmp_2_cfg_a,
  input         io_pmp_2_cfg_x,
  input         io_pmp_2_cfg_w,
  input         io_pmp_2_cfg_r,
  input  [29:0] io_pmp_2_addr,
  input  [31:0] io_pmp_2_mask,
  input         io_pmp_3_cfg_l,
  input  [1:0]  io_pmp_3_cfg_a,
  input         io_pmp_3_cfg_x,
  input         io_pmp_3_cfg_w,
  input         io_pmp_3_cfg_r,
  input  [29:0] io_pmp_3_addr,
  input  [31:0] io_pmp_3_mask,
  input         io_pmp_4_cfg_l,
  input  [1:0]  io_pmp_4_cfg_a,
  input         io_pmp_4_cfg_x,
  input         io_pmp_4_cfg_w,
  input         io_pmp_4_cfg_r,
  input  [29:0] io_pmp_4_addr,
  input  [31:0] io_pmp_4_mask,
  input         io_pmp_5_cfg_l,
  input  [1:0]  io_pmp_5_cfg_a,
  input         io_pmp_5_cfg_x,
  input         io_pmp_5_cfg_w,
  input         io_pmp_5_cfg_r,
  input  [29:0] io_pmp_5_addr,
  input  [31:0] io_pmp_5_mask,
  input         io_pmp_6_cfg_l,
  input  [1:0]  io_pmp_6_cfg_a,
  input         io_pmp_6_cfg_x,
  input         io_pmp_6_cfg_w,
  input         io_pmp_6_cfg_r,
  input  [29:0] io_pmp_6_addr,
  input  [31:0] io_pmp_6_mask,
  input         io_pmp_7_cfg_l,
  input  [1:0]  io_pmp_7_cfg_a,
  input         io_pmp_7_cfg_x,
  input         io_pmp_7_cfg_w,
  input         io_pmp_7_cfg_r,
  input  [29:0] io_pmp_7_addr,
  input  [31:0] io_pmp_7_mask,
  input  [31:0] io_addr,
  output        io_r,
  output        io_w,
  output        io_x,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  default_; // @[PMP.scala 157:56]
  wire [31:0] _T_2; // @[PMP.scala 62:36]
  wire [31:0] _T_4; // @[PMP.scala 62:48]
  wire [31:0] _T_6; // @[PMP.scala 65:47]
  wire [31:0] _T_8; // @[PMP.scala 65:52]
  wire  _T_9; // @[PMP.scala 65:58]
  wire [31:0] _T_15; // @[PMP.scala 62:36]
  wire [31:0] _T_17; // @[PMP.scala 62:48]
  wire  _T_19; // @[PMP.scala 79:9]
  wire  _T_25; // @[PMP.scala 79:9]
  wire  _T_26; // @[PMP.scala 96:48]
  wire  _T_27; // @[PMP.scala 134:61]
  wire  _T_28; // @[PMP.scala 134:8]
  wire  _T_30; // @[PMP.scala 165:26]
  wire  _T_82; // @[PMP.scala 183:40]
  wire  _T_84; // @[PMP.scala 184:40]
  wire  _T_86; // @[PMP.scala 185:40]
  wire  _T_88_cfg_x; // @[PMP.scala 186:8]
  wire  _T_88_cfg_w; // @[PMP.scala 186:8]
  wire  _T_88_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_94; // @[PMP.scala 65:47]
  wire [31:0] _T_96; // @[PMP.scala 65:52]
  wire  _T_97; // @[PMP.scala 65:58]
  wire [31:0] _T_103; // @[PMP.scala 62:36]
  wire [31:0] _T_105; // @[PMP.scala 62:48]
  wire  _T_107; // @[PMP.scala 79:9]
  wire  _T_114; // @[PMP.scala 96:48]
  wire  _T_115; // @[PMP.scala 134:61]
  wire  _T_116; // @[PMP.scala 134:8]
  wire  _T_118; // @[PMP.scala 165:26]
  wire  _T_170; // @[PMP.scala 183:40]
  wire  _T_172; // @[PMP.scala 184:40]
  wire  _T_174; // @[PMP.scala 185:40]
  wire  _T_176_cfg_x; // @[PMP.scala 186:8]
  wire  _T_176_cfg_w; // @[PMP.scala 186:8]
  wire  _T_176_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_182; // @[PMP.scala 65:47]
  wire [31:0] _T_184; // @[PMP.scala 65:52]
  wire  _T_185; // @[PMP.scala 65:58]
  wire [31:0] _T_191; // @[PMP.scala 62:36]
  wire [31:0] _T_193; // @[PMP.scala 62:48]
  wire  _T_195; // @[PMP.scala 79:9]
  wire  _T_202; // @[PMP.scala 96:48]
  wire  _T_203; // @[PMP.scala 134:61]
  wire  _T_204; // @[PMP.scala 134:8]
  wire  _T_206; // @[PMP.scala 165:26]
  wire  _T_258; // @[PMP.scala 183:40]
  wire  _T_260; // @[PMP.scala 184:40]
  wire  _T_262; // @[PMP.scala 185:40]
  wire  _T_264_cfg_x; // @[PMP.scala 186:8]
  wire  _T_264_cfg_w; // @[PMP.scala 186:8]
  wire  _T_264_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_270; // @[PMP.scala 65:47]
  wire [31:0] _T_272; // @[PMP.scala 65:52]
  wire  _T_273; // @[PMP.scala 65:58]
  wire [31:0] _T_279; // @[PMP.scala 62:36]
  wire [31:0] _T_281; // @[PMP.scala 62:48]
  wire  _T_283; // @[PMP.scala 79:9]
  wire  _T_290; // @[PMP.scala 96:48]
  wire  _T_291; // @[PMP.scala 134:61]
  wire  _T_292; // @[PMP.scala 134:8]
  wire  _T_294; // @[PMP.scala 165:26]
  wire  _T_346; // @[PMP.scala 183:40]
  wire  _T_348; // @[PMP.scala 184:40]
  wire  _T_350; // @[PMP.scala 185:40]
  wire  _T_352_cfg_x; // @[PMP.scala 186:8]
  wire  _T_352_cfg_w; // @[PMP.scala 186:8]
  wire  _T_352_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_358; // @[PMP.scala 65:47]
  wire [31:0] _T_360; // @[PMP.scala 65:52]
  wire  _T_361; // @[PMP.scala 65:58]
  wire [31:0] _T_367; // @[PMP.scala 62:36]
  wire [31:0] _T_369; // @[PMP.scala 62:48]
  wire  _T_371; // @[PMP.scala 79:9]
  wire  _T_378; // @[PMP.scala 96:48]
  wire  _T_379; // @[PMP.scala 134:61]
  wire  _T_380; // @[PMP.scala 134:8]
  wire  _T_382; // @[PMP.scala 165:26]
  wire  _T_434; // @[PMP.scala 183:40]
  wire  _T_436; // @[PMP.scala 184:40]
  wire  _T_438; // @[PMP.scala 185:40]
  wire  _T_440_cfg_x; // @[PMP.scala 186:8]
  wire  _T_440_cfg_w; // @[PMP.scala 186:8]
  wire  _T_440_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_446; // @[PMP.scala 65:47]
  wire [31:0] _T_448; // @[PMP.scala 65:52]
  wire  _T_449; // @[PMP.scala 65:58]
  wire [31:0] _T_455; // @[PMP.scala 62:36]
  wire [31:0] _T_457; // @[PMP.scala 62:48]
  wire  _T_459; // @[PMP.scala 79:9]
  wire  _T_466; // @[PMP.scala 96:48]
  wire  _T_467; // @[PMP.scala 134:61]
  wire  _T_468; // @[PMP.scala 134:8]
  wire  _T_470; // @[PMP.scala 165:26]
  wire  _T_522; // @[PMP.scala 183:40]
  wire  _T_524; // @[PMP.scala 184:40]
  wire  _T_526; // @[PMP.scala 185:40]
  wire  _T_528_cfg_x; // @[PMP.scala 186:8]
  wire  _T_528_cfg_w; // @[PMP.scala 186:8]
  wire  _T_528_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_534; // @[PMP.scala 65:47]
  wire [31:0] _T_536; // @[PMP.scala 65:52]
  wire  _T_537; // @[PMP.scala 65:58]
  wire [31:0] _T_543; // @[PMP.scala 62:36]
  wire [31:0] _T_545; // @[PMP.scala 62:48]
  wire  _T_547; // @[PMP.scala 79:9]
  wire  _T_554; // @[PMP.scala 96:48]
  wire  _T_555; // @[PMP.scala 134:61]
  wire  _T_556; // @[PMP.scala 134:8]
  wire  _T_558; // @[PMP.scala 165:26]
  wire  _T_610; // @[PMP.scala 183:40]
  wire  _T_612; // @[PMP.scala 184:40]
  wire  _T_614; // @[PMP.scala 185:40]
  wire  _T_616_cfg_x; // @[PMP.scala 186:8]
  wire  _T_616_cfg_w; // @[PMP.scala 186:8]
  wire  _T_616_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_622; // @[PMP.scala 65:47]
  wire [31:0] _T_624; // @[PMP.scala 65:52]
  wire  _T_625; // @[PMP.scala 65:58]
  wire  _T_643; // @[PMP.scala 134:61]
  wire  _T_644; // @[PMP.scala 134:8]
  wire  _T_646; // @[PMP.scala 165:26]
  wire  _T_698; // @[PMP.scala 183:40]
  wire  _T_700; // @[PMP.scala 184:40]
  wire  _T_702; // @[PMP.scala 185:40]
  wire [29:0] PMPChecker_2_covSum;
  assign default_ = io_prv > 2'h1; // @[PMP.scala 157:56]
  assign _T_2 = {io_pmp_7_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_4 = ~_T_2 | 32'h3; // @[PMP.scala 62:48]
  assign _T_6 = io_addr ^ ~_T_4; // @[PMP.scala 65:47]
  assign _T_8 = _T_6 & ~io_pmp_7_mask; // @[PMP.scala 65:52]
  assign _T_9 = _T_8 == 32'h0; // @[PMP.scala 65:58]
  assign _T_15 = {io_pmp_6_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_17 = ~_T_15 | 32'h3; // @[PMP.scala 62:48]
  assign _T_19 = io_addr < ~_T_17; // @[PMP.scala 79:9]
  assign _T_25 = io_addr < ~_T_4; // @[PMP.scala 79:9]
  assign _T_26 = ~_T_19 & _T_25; // @[PMP.scala 96:48]
  assign _T_27 = io_pmp_7_cfg_a[0] & _T_26; // @[PMP.scala 134:61]
  assign _T_28 = io_pmp_7_cfg_a[1] ? _T_9 : _T_27; // @[PMP.scala 134:8]
  assign _T_30 = default_ & ~io_pmp_7_cfg_l; // @[PMP.scala 165:26]
  assign _T_82 = io_pmp_7_cfg_r | _T_30; // @[PMP.scala 183:40]
  assign _T_84 = io_pmp_7_cfg_w | _T_30; // @[PMP.scala 184:40]
  assign _T_86 = io_pmp_7_cfg_x | _T_30; // @[PMP.scala 185:40]
  assign _T_88_cfg_x = _T_28 ? _T_86 : default_; // @[PMP.scala 186:8]
  assign _T_88_cfg_w = _T_28 ? _T_84 : default_; // @[PMP.scala 186:8]
  assign _T_88_cfg_r = _T_28 ? _T_82 : default_; // @[PMP.scala 186:8]
  assign _T_94 = io_addr ^ ~_T_17; // @[PMP.scala 65:47]
  assign _T_96 = _T_94 & ~io_pmp_6_mask; // @[PMP.scala 65:52]
  assign _T_97 = _T_96 == 32'h0; // @[PMP.scala 65:58]
  assign _T_103 = {io_pmp_5_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_105 = ~_T_103 | 32'h3; // @[PMP.scala 62:48]
  assign _T_107 = io_addr < ~_T_105; // @[PMP.scala 79:9]
  assign _T_114 = ~_T_107 & _T_19; // @[PMP.scala 96:48]
  assign _T_115 = io_pmp_6_cfg_a[0] & _T_114; // @[PMP.scala 134:61]
  assign _T_116 = io_pmp_6_cfg_a[1] ? _T_97 : _T_115; // @[PMP.scala 134:8]
  assign _T_118 = default_ & ~io_pmp_6_cfg_l; // @[PMP.scala 165:26]
  assign _T_170 = io_pmp_6_cfg_r | _T_118; // @[PMP.scala 183:40]
  assign _T_172 = io_pmp_6_cfg_w | _T_118; // @[PMP.scala 184:40]
  assign _T_174 = io_pmp_6_cfg_x | _T_118; // @[PMP.scala 185:40]
  assign _T_176_cfg_x = _T_116 ? _T_174 : _T_88_cfg_x; // @[PMP.scala 186:8]
  assign _T_176_cfg_w = _T_116 ? _T_172 : _T_88_cfg_w; // @[PMP.scala 186:8]
  assign _T_176_cfg_r = _T_116 ? _T_170 : _T_88_cfg_r; // @[PMP.scala 186:8]
  assign _T_182 = io_addr ^ ~_T_105; // @[PMP.scala 65:47]
  assign _T_184 = _T_182 & ~io_pmp_5_mask; // @[PMP.scala 65:52]
  assign _T_185 = _T_184 == 32'h0; // @[PMP.scala 65:58]
  assign _T_191 = {io_pmp_4_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_193 = ~_T_191 | 32'h3; // @[PMP.scala 62:48]
  assign _T_195 = io_addr < ~_T_193; // @[PMP.scala 79:9]
  assign _T_202 = ~_T_195 & _T_107; // @[PMP.scala 96:48]
  assign _T_203 = io_pmp_5_cfg_a[0] & _T_202; // @[PMP.scala 134:61]
  assign _T_204 = io_pmp_5_cfg_a[1] ? _T_185 : _T_203; // @[PMP.scala 134:8]
  assign _T_206 = default_ & ~io_pmp_5_cfg_l; // @[PMP.scala 165:26]
  assign _T_258 = io_pmp_5_cfg_r | _T_206; // @[PMP.scala 183:40]
  assign _T_260 = io_pmp_5_cfg_w | _T_206; // @[PMP.scala 184:40]
  assign _T_262 = io_pmp_5_cfg_x | _T_206; // @[PMP.scala 185:40]
  assign _T_264_cfg_x = _T_204 ? _T_262 : _T_176_cfg_x; // @[PMP.scala 186:8]
  assign _T_264_cfg_w = _T_204 ? _T_260 : _T_176_cfg_w; // @[PMP.scala 186:8]
  assign _T_264_cfg_r = _T_204 ? _T_258 : _T_176_cfg_r; // @[PMP.scala 186:8]
  assign _T_270 = io_addr ^ ~_T_193; // @[PMP.scala 65:47]
  assign _T_272 = _T_270 & ~io_pmp_4_mask; // @[PMP.scala 65:52]
  assign _T_273 = _T_272 == 32'h0; // @[PMP.scala 65:58]
  assign _T_279 = {io_pmp_3_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_281 = ~_T_279 | 32'h3; // @[PMP.scala 62:48]
  assign _T_283 = io_addr < ~_T_281; // @[PMP.scala 79:9]
  assign _T_290 = ~_T_283 & _T_195; // @[PMP.scala 96:48]
  assign _T_291 = io_pmp_4_cfg_a[0] & _T_290; // @[PMP.scala 134:61]
  assign _T_292 = io_pmp_4_cfg_a[1] ? _T_273 : _T_291; // @[PMP.scala 134:8]
  assign _T_294 = default_ & ~io_pmp_4_cfg_l; // @[PMP.scala 165:26]
  assign _T_346 = io_pmp_4_cfg_r | _T_294; // @[PMP.scala 183:40]
  assign _T_348 = io_pmp_4_cfg_w | _T_294; // @[PMP.scala 184:40]
  assign _T_350 = io_pmp_4_cfg_x | _T_294; // @[PMP.scala 185:40]
  assign _T_352_cfg_x = _T_292 ? _T_350 : _T_264_cfg_x; // @[PMP.scala 186:8]
  assign _T_352_cfg_w = _T_292 ? _T_348 : _T_264_cfg_w; // @[PMP.scala 186:8]
  assign _T_352_cfg_r = _T_292 ? _T_346 : _T_264_cfg_r; // @[PMP.scala 186:8]
  assign _T_358 = io_addr ^ ~_T_281; // @[PMP.scala 65:47]
  assign _T_360 = _T_358 & ~io_pmp_3_mask; // @[PMP.scala 65:52]
  assign _T_361 = _T_360 == 32'h0; // @[PMP.scala 65:58]
  assign _T_367 = {io_pmp_2_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_369 = ~_T_367 | 32'h3; // @[PMP.scala 62:48]
  assign _T_371 = io_addr < ~_T_369; // @[PMP.scala 79:9]
  assign _T_378 = ~_T_371 & _T_283; // @[PMP.scala 96:48]
  assign _T_379 = io_pmp_3_cfg_a[0] & _T_378; // @[PMP.scala 134:61]
  assign _T_380 = io_pmp_3_cfg_a[1] ? _T_361 : _T_379; // @[PMP.scala 134:8]
  assign _T_382 = default_ & ~io_pmp_3_cfg_l; // @[PMP.scala 165:26]
  assign _T_434 = io_pmp_3_cfg_r | _T_382; // @[PMP.scala 183:40]
  assign _T_436 = io_pmp_3_cfg_w | _T_382; // @[PMP.scala 184:40]
  assign _T_438 = io_pmp_3_cfg_x | _T_382; // @[PMP.scala 185:40]
  assign _T_440_cfg_x = _T_380 ? _T_438 : _T_352_cfg_x; // @[PMP.scala 186:8]
  assign _T_440_cfg_w = _T_380 ? _T_436 : _T_352_cfg_w; // @[PMP.scala 186:8]
  assign _T_440_cfg_r = _T_380 ? _T_434 : _T_352_cfg_r; // @[PMP.scala 186:8]
  assign _T_446 = io_addr ^ ~_T_369; // @[PMP.scala 65:47]
  assign _T_448 = _T_446 & ~io_pmp_2_mask; // @[PMP.scala 65:52]
  assign _T_449 = _T_448 == 32'h0; // @[PMP.scala 65:58]
  assign _T_455 = {io_pmp_1_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_457 = ~_T_455 | 32'h3; // @[PMP.scala 62:48]
  assign _T_459 = io_addr < ~_T_457; // @[PMP.scala 79:9]
  assign _T_466 = ~_T_459 & _T_371; // @[PMP.scala 96:48]
  assign _T_467 = io_pmp_2_cfg_a[0] & _T_466; // @[PMP.scala 134:61]
  assign _T_468 = io_pmp_2_cfg_a[1] ? _T_449 : _T_467; // @[PMP.scala 134:8]
  assign _T_470 = default_ & ~io_pmp_2_cfg_l; // @[PMP.scala 165:26]
  assign _T_522 = io_pmp_2_cfg_r | _T_470; // @[PMP.scala 183:40]
  assign _T_524 = io_pmp_2_cfg_w | _T_470; // @[PMP.scala 184:40]
  assign _T_526 = io_pmp_2_cfg_x | _T_470; // @[PMP.scala 185:40]
  assign _T_528_cfg_x = _T_468 ? _T_526 : _T_440_cfg_x; // @[PMP.scala 186:8]
  assign _T_528_cfg_w = _T_468 ? _T_524 : _T_440_cfg_w; // @[PMP.scala 186:8]
  assign _T_528_cfg_r = _T_468 ? _T_522 : _T_440_cfg_r; // @[PMP.scala 186:8]
  assign _T_534 = io_addr ^ ~_T_457; // @[PMP.scala 65:47]
  assign _T_536 = _T_534 & ~io_pmp_1_mask; // @[PMP.scala 65:52]
  assign _T_537 = _T_536 == 32'h0; // @[PMP.scala 65:58]
  assign _T_543 = {io_pmp_0_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _T_545 = ~_T_543 | 32'h3; // @[PMP.scala 62:48]
  assign _T_547 = io_addr < ~_T_545; // @[PMP.scala 79:9]
  assign _T_554 = ~_T_547 & _T_459; // @[PMP.scala 96:48]
  assign _T_555 = io_pmp_1_cfg_a[0] & _T_554; // @[PMP.scala 134:61]
  assign _T_556 = io_pmp_1_cfg_a[1] ? _T_537 : _T_555; // @[PMP.scala 134:8]
  assign _T_558 = default_ & ~io_pmp_1_cfg_l; // @[PMP.scala 165:26]
  assign _T_610 = io_pmp_1_cfg_r | _T_558; // @[PMP.scala 183:40]
  assign _T_612 = io_pmp_1_cfg_w | _T_558; // @[PMP.scala 184:40]
  assign _T_614 = io_pmp_1_cfg_x | _T_558; // @[PMP.scala 185:40]
  assign _T_616_cfg_x = _T_556 ? _T_614 : _T_528_cfg_x; // @[PMP.scala 186:8]
  assign _T_616_cfg_w = _T_556 ? _T_612 : _T_528_cfg_w; // @[PMP.scala 186:8]
  assign _T_616_cfg_r = _T_556 ? _T_610 : _T_528_cfg_r; // @[PMP.scala 186:8]
  assign _T_622 = io_addr ^ ~_T_545; // @[PMP.scala 65:47]
  assign _T_624 = _T_622 & ~io_pmp_0_mask; // @[PMP.scala 65:52]
  assign _T_625 = _T_624 == 32'h0; // @[PMP.scala 65:58]
  assign _T_643 = io_pmp_0_cfg_a[0] & _T_547; // @[PMP.scala 134:61]
  assign _T_644 = io_pmp_0_cfg_a[1] ? _T_625 : _T_643; // @[PMP.scala 134:8]
  assign _T_646 = default_ & ~io_pmp_0_cfg_l; // @[PMP.scala 165:26]
  assign _T_698 = io_pmp_0_cfg_r | _T_646; // @[PMP.scala 183:40]
  assign _T_700 = io_pmp_0_cfg_w | _T_646; // @[PMP.scala 184:40]
  assign _T_702 = io_pmp_0_cfg_x | _T_646; // @[PMP.scala 185:40]
  assign io_r = _T_644 ? _T_698 : _T_616_cfg_r; // @[PMP.scala 189:8]
  assign io_w = _T_644 ? _T_700 : _T_616_cfg_w; // @[PMP.scala 190:8]
  assign io_x = _T_644 ? _T_702 : _T_616_cfg_x; // @[PMP.scala 191:8]
  assign PMPChecker_2_covSum = 30'h0;
  assign io_covSum = PMPChecker_2_covSum;
  assign metaAssert = 1'h0;
endmodule
module NonSyncResetSynchronizerPrimitiveShiftReg_d3(
  input         clock,
  input         io_d,
  output        io_q,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  sync_0; // @[SynchronizerReg.scala 59:68]
  reg [31:0] _RAND_0;
  reg  sync_1; // @[SynchronizerReg.scala 59:68]
  reg [31:0] _RAND_1;
  reg  sync_2; // @[SynchronizerReg.scala 59:68]
  reg [31:0] _RAND_2;
  wire [29:0] NonSyncResetSynchronizerPrimitiveShiftReg_d3_covSum;
  assign io_q = sync_0; // @[SynchronizerReg.scala 67:10]
  assign NonSyncResetSynchronizerPrimitiveShiftReg_d3_covSum = 30'h0;
  assign io_covSum = NonSyncResetSynchronizerPrimitiveShiftReg_d3_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sync_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sync_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  sync_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      sync_0 <= 1'h0;
    end else begin
      sync_0 <= sync_1;
    end
    if (metaReset) begin
      sync_1 <= 1'h0;
    end else begin
      sync_1 <= sync_2;
    end
    if (metaReset) begin
      sync_2 <= 1'h0;
    end else begin
      sync_2 <= io_d;
    end
  end
endmodule
module MulAddRecFNPipe(
  input         clock,
  input         reset,
  input         io_validin,
  input  [1:0]  io_op,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [1:0] mulAddRecFNToRaw_preMul_io_op; // @[FPU.scala 600:41]
  wire [32:0] mulAddRecFNToRaw_preMul_io_a; // @[FPU.scala 600:41]
  wire [32:0] mulAddRecFNToRaw_preMul_io_b; // @[FPU.scala 600:41]
  wire [32:0] mulAddRecFNToRaw_preMul_io_c; // @[FPU.scala 600:41]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[FPU.scala 600:41]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[FPU.scala 600:41]
  wire [47:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FPU.scala 600:41]
  wire [9:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FPU.scala 600:41]
  wire [4:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FPU.scala 600:41]
  wire [25:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FPU.scala 600:41]
  wire [29:0] mulAddRecFNToRaw_preMul_io_covSum; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_metaAssert; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[FPU.scala 601:42]
  wire [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[FPU.scala 601:42]
  wire [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[FPU.scala 601:42]
  wire [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[FPU.scala 601:42]
  wire [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[FPU.scala 601:42]
  wire [2:0] mulAddRecFNToRaw_postMul_io_roundingMode; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FPU.scala 601:42]
  wire [9:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FPU.scala 601:42]
  wire [26:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FPU.scala 601:42]
  wire [29:0] mulAddRecFNToRaw_postMul_io_covSum; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_metaAssert; // @[FPU.scala 601:42]
  wire  roundRawFNToRecFN_io_invalidExc; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_io_in_isInf; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_io_in_isZero; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_io_in_sign; // @[FPU.scala 628:35]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[FPU.scala 628:35]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[FPU.scala 628:35]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_io_detectTininess; // @[FPU.scala 628:35]
  wire [32:0] roundRawFNToRecFN_io_out; // @[FPU.scala 628:35]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[FPU.scala 628:35]
  wire [29:0] roundRawFNToRecFN_io_covSum; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_metaAssert; // @[FPU.scala 628:35]
  wire [47:0] _T; // @[FPU.scala 609:45]
  wire [48:0] mulAddResult; // @[FPU.scala 610:50]
  reg  _T_2_isSigNaNAny; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg  _T_2_isNaNAOrB; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  _T_2_isInfA; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg  _T_2_isZeroA; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg  _T_2_isInfB; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  _T_2_isZeroB; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  _T_2_signProd; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  _T_2_isNaNC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg  _T_2_isInfC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg  _T_2_isZeroC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [9:0] _T_2_sExpSum; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg  _T_2_doSubMags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg  _T_2_CIsDominant; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [4:0] _T_2_CDom_CAlignDist; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [25:0] _T_2_highAlignedSigC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg  _T_2_bit0AlignedSigC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [48:0] _T_5; // @[Reg.scala 15:16]
  reg [63:0] _RAND_16;
  reg [2:0] _T_8; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [2:0] roundingMode_stage0; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg  detectTininess_stage0; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg  valid_stage0; // @[Valid.scala 117:22]
  reg [31:0] _RAND_20;
  reg  _T_20; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg  _T_23_isNaN; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg  _T_23_isInf; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg  _T_23_isZero; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg  _T_23_sign; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [9:0] _T_23_sExp; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [26:0] _T_23_sig; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [2:0] _T_26; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg  _T_29; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg  MulAddRecFNPipe_state; // @[Register tracking MulAddRecFNPipe state]
  reg [31:0] _RAND_30;
  reg  MulAddRecFNPipe_cov [0:1]; // @[Coverage map for MulAddRecFNPipe]
  reg [31:0] _RAND_31;
  wire  MulAddRecFNPipe_cov_read_data; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_read_addr; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_write_data; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_write_addr; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_write_mask; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_write_en; // @[Coverage map for MulAddRecFNPipe]
  reg [29:0] MulAddRecFNPipe_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_32;
  wire  valid_stage0_shl;
  wire  valid_stage0_pad;
  wire [29:0] mulAddRecFNToRaw_preMul_sum;
  wire [29:0] mulAddRecFNToRaw_postMul_sum;
  wire [29:0] roundRawFNToRecFN_sum;
  wire  mulAddRecFNToRaw_preMul_metaAssert_wire;
  wire  mulAddRecFNToRaw_postMul_metaAssert_wire;
  wire  roundRawFNToRecFN_metaAssert_wire;
  wire  MulAddRecFNPipe_or2;
  wire  MulAddRecFNPipe_or0;
  reg  MulAddRecFNPipe_metaAssert;
  reg [31:0] _RAND_33;
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[FPU.scala 600:41]
    .io_op(mulAddRecFNToRaw_preMul_io_op),
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC),
    .io_covSum(mulAddRecFNToRaw_preMul_io_covSum),
    .metaAssert(mulAddRecFNToRaw_preMul_metaAssert)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[FPU.scala 601:42]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_roundingMode(mulAddRecFNToRaw_postMul_io_roundingMode),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig),
    .io_covSum(mulAddRecFNToRaw_postMul_io_covSum),
    .metaAssert(mulAddRecFNToRaw_postMul_metaAssert)
  );
  RoundRawFNToRecFN_2 roundRawFNToRecFN ( // @[FPU.scala 628:35]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundRawFNToRecFN_io_covSum),
    .metaAssert(roundRawFNToRecFN_metaAssert)
  );
  assign _T = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB; // @[FPU.scala 609:45]
  assign mulAddResult = _T + mulAddRecFNToRaw_preMul_io_mulAddC; // @[FPU.scala 610:50]
  assign io_out = roundRawFNToRecFN_io_out; // @[FPU.scala 639:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[FPU.scala 640:23]
  assign mulAddRecFNToRaw_preMul_io_op = io_op; // @[FPU.scala 603:35]
  assign mulAddRecFNToRaw_preMul_io_a = io_a; // @[FPU.scala 604:35]
  assign mulAddRecFNToRaw_preMul_io_b = io_b; // @[FPU.scala 605:35]
  assign mulAddRecFNToRaw_preMul_io_c = io_c; // @[FPU.scala 606:35]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = _T_2_isSigNaNAny; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = _T_2_isNaNAOrB; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = _T_2_isInfA; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = _T_2_isZeroA; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = _T_2_isInfB; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = _T_2_isZeroB; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = _T_2_signProd; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = _T_2_isNaNC; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = _T_2_isInfC; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = _T_2_isZeroC; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = _T_2_sExpSum; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = _T_2_doSubMags; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = _T_2_CIsDominant; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = _T_2_CDom_CAlignDist; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = _T_2_highAlignedSigC; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = _T_2_bit0AlignedSigC; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T_5; // @[FPU.scala 619:46]
  assign mulAddRecFNToRaw_postMul_io_roundingMode = _T_8; // @[FPU.scala 620:46]
  assign roundRawFNToRecFN_io_invalidExc = _T_20; // @[FPU.scala 631:45]
  assign roundRawFNToRecFN_io_infiniteExc = 1'h0; // @[FPU.scala 637:38]
  assign roundRawFNToRecFN_io_in_isNaN = _T_23_isNaN; // @[FPU.scala 632:45]
  assign roundRawFNToRecFN_io_in_isInf = _T_23_isInf; // @[FPU.scala 632:45]
  assign roundRawFNToRecFN_io_in_isZero = _T_23_isZero; // @[FPU.scala 632:45]
  assign roundRawFNToRecFN_io_in_sign = _T_23_sign; // @[FPU.scala 632:45]
  assign roundRawFNToRecFN_io_in_sExp = _T_23_sExp; // @[FPU.scala 632:45]
  assign roundRawFNToRecFN_io_in_sig = _T_23_sig; // @[FPU.scala 632:45]
  assign roundRawFNToRecFN_io_roundingMode = _T_26; // @[FPU.scala 633:45]
  assign roundRawFNToRecFN_io_detectTininess = _T_29; // @[FPU.scala 634:45]
  assign MulAddRecFNPipe_cov_read_addr = MulAddRecFNPipe_state;
  assign MulAddRecFNPipe_cov_read_data = MulAddRecFNPipe_cov[MulAddRecFNPipe_cov_read_addr]; // @[Coverage map for MulAddRecFNPipe]
  assign MulAddRecFNPipe_cov_write_data = 1'h1;
  assign MulAddRecFNPipe_cov_write_addr = MulAddRecFNPipe_state;
  assign MulAddRecFNPipe_cov_write_mask = 1'h1;
  assign MulAddRecFNPipe_cov_write_en = 1'h1;
  assign valid_stage0_shl = valid_stage0;
  assign valid_stage0_pad = valid_stage0_shl;
  assign mulAddRecFNToRaw_preMul_sum = MulAddRecFNPipe_covSum + mulAddRecFNToRaw_preMul_io_covSum;
  assign mulAddRecFNToRaw_postMul_sum = mulAddRecFNToRaw_preMul_sum + mulAddRecFNToRaw_postMul_io_covSum;
  assign roundRawFNToRecFN_sum = mulAddRecFNToRaw_postMul_sum + roundRawFNToRecFN_io_covSum;
  assign io_covSum = roundRawFNToRecFN_sum;
  assign mulAddRecFNToRaw_preMul_metaAssert_wire = mulAddRecFNToRaw_preMul_metaAssert;
  assign mulAddRecFNToRaw_postMul_metaAssert_wire = mulAddRecFNToRaw_postMul_metaAssert;
  assign roundRawFNToRecFN_metaAssert_wire = roundRawFNToRecFN_metaAssert;
  assign MulAddRecFNPipe_or2 = mulAddRecFNToRaw_postMul_metaAssert_wire | roundRawFNToRecFN_metaAssert_wire;
  assign MulAddRecFNPipe_or0 = mulAddRecFNToRaw_preMul_metaAssert_wire | MulAddRecFNPipe_or2;
  assign metaAssert = MulAddRecFNPipe_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2_isSigNaNAny = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2_isNaNAOrB = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_isInfA = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2_isZeroA = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2_isInfB = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2_isZeroB = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2_signProd = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2_isNaNC = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2_isInfC = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_2_isZeroC = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2_sExpSum = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2_doSubMags = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2_CIsDominant = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2_CDom_CAlignDist = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_2_highAlignedSigC = _RAND_14[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2_bit0AlignedSigC = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  _T_5 = _RAND_16[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_8 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  roundingMode_stage0 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  detectTininess_stage0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  valid_stage0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_20 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_23_isNaN = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_23_isInf = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_23_isZero = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_23_sign = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_23_sExp = _RAND_26[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_23_sig = _RAND_27[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_26 = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  MulAddRecFNPipe_state = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    MulAddRecFNPipe_cov[initvar] = _RAND_31[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  MulAddRecFNPipe_covSum = _RAND_32[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  MulAddRecFNPipe_metaAssert = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_2_isSigNaNAny <= 1'h0;
    end else if (io_validin) begin
      _T_2_isSigNaNAny <= mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny;
    end
    if (metaReset) begin
      _T_2_isNaNAOrB <= 1'h0;
    end else if (io_validin) begin
      _T_2_isNaNAOrB <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB;
    end
    if (metaReset) begin
      _T_2_isInfA <= 1'h0;
    end else if (io_validin) begin
      _T_2_isInfA <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfA;
    end
    if (metaReset) begin
      _T_2_isZeroA <= 1'h0;
    end else if (io_validin) begin
      _T_2_isZeroA <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA;
    end
    if (metaReset) begin
      _T_2_isInfB <= 1'h0;
    end else if (io_validin) begin
      _T_2_isInfB <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfB;
    end
    if (metaReset) begin
      _T_2_isZeroB <= 1'h0;
    end else if (io_validin) begin
      _T_2_isZeroB <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB;
    end
    if (metaReset) begin
      _T_2_signProd <= 1'h0;
    end else if (io_validin) begin
      _T_2_signProd <= mulAddRecFNToRaw_preMul_io_toPostMul_signProd;
    end
    if (metaReset) begin
      _T_2_isNaNC <= 1'h0;
    end else if (io_validin) begin
      _T_2_isNaNC <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC;
    end
    if (metaReset) begin
      _T_2_isInfC <= 1'h0;
    end else if (io_validin) begin
      _T_2_isInfC <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfC;
    end
    if (metaReset) begin
      _T_2_isZeroC <= 1'h0;
    end else if (io_validin) begin
      _T_2_isZeroC <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC;
    end
    if (metaReset) begin
      _T_2_sExpSum <= 10'h0;
    end else if (io_validin) begin
      _T_2_sExpSum <= mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum;
    end
    if (metaReset) begin
      _T_2_doSubMags <= 1'h0;
    end else if (io_validin) begin
      _T_2_doSubMags <= mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags;
    end
    if (metaReset) begin
      _T_2_CIsDominant <= 1'h0;
    end else if (io_validin) begin
      _T_2_CIsDominant <= mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant;
    end
    if (metaReset) begin
      _T_2_CDom_CAlignDist <= 5'h0;
    end else if (io_validin) begin
      _T_2_CDom_CAlignDist <= mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist;
    end
    if (metaReset) begin
      _T_2_highAlignedSigC <= 26'h0;
    end else if (io_validin) begin
      _T_2_highAlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC;
    end
    if (metaReset) begin
      _T_2_bit0AlignedSigC <= 1'h0;
    end else if (io_validin) begin
      _T_2_bit0AlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC;
    end
    if (metaReset) begin
      _T_5 <= 49'h0;
    end else if (io_validin) begin
      _T_5 <= mulAddResult;
    end
    if (metaReset) begin
      _T_8 <= 3'h0;
    end else if (io_validin) begin
      _T_8 <= io_roundingMode;
    end
    if (metaReset) begin
      roundingMode_stage0 <= 3'h0;
    end else if (io_validin) begin
      roundingMode_stage0 <= io_roundingMode;
    end
    if (metaReset) begin
      detectTininess_stage0 <= 1'h0;
    end else begin
      detectTininess_stage0 <= io_validin | detectTininess_stage0;
    end
    if (metaReset) begin
      valid_stage0 <= 1'h0;
    end else if (reset) begin
      valid_stage0 <= 1'h0;
    end else begin
      valid_stage0 <= io_validin;
    end
    if (metaReset) begin
      _T_20 <= 1'h0;
    end else if (valid_stage0) begin
      _T_20 <= mulAddRecFNToRaw_postMul_io_invalidExc;
    end
    if (metaReset) begin
      _T_23_isNaN <= 1'h0;
    end else if (valid_stage0) begin
      _T_23_isNaN <= mulAddRecFNToRaw_postMul_io_rawOut_isNaN;
    end
    if (metaReset) begin
      _T_23_isInf <= 1'h0;
    end else if (valid_stage0) begin
      _T_23_isInf <= mulAddRecFNToRaw_postMul_io_rawOut_isInf;
    end
    if (metaReset) begin
      _T_23_isZero <= 1'h0;
    end else if (valid_stage0) begin
      _T_23_isZero <= mulAddRecFNToRaw_postMul_io_rawOut_isZero;
    end
    if (metaReset) begin
      _T_23_sign <= 1'h0;
    end else if (valid_stage0) begin
      _T_23_sign <= mulAddRecFNToRaw_postMul_io_rawOut_sign;
    end
    if (metaReset) begin
      _T_23_sExp <= 10'h0;
    end else if (valid_stage0) begin
      _T_23_sExp <= mulAddRecFNToRaw_postMul_io_rawOut_sExp;
    end
    if (metaReset) begin
      _T_23_sig <= 27'h0;
    end else if (valid_stage0) begin
      _T_23_sig <= mulAddRecFNToRaw_postMul_io_rawOut_sig;
    end
    if (metaReset) begin
      _T_26 <= 3'h0;
    end else if (valid_stage0) begin
      _T_26 <= roundingMode_stage0;
    end
    if (metaReset) begin
      _T_29 <= 1'h0;
    end else if (valid_stage0) begin
      _T_29 <= detectTininess_stage0;
    end
    MulAddRecFNPipe_state <= valid_stage0_pad;
    if (!(MulAddRecFNPipe_cov_read_data)) begin
      MulAddRecFNPipe_covSum <= MulAddRecFNPipe_covSum + 1'h1;
    end
    if (metaReset) begin
      MulAddRecFNPipe_metaAssert <= 1'h0;
    end else begin
      MulAddRecFNPipe_metaAssert <= MulAddRecFNPipe_metaAssert | MulAddRecFNPipe_or0;
    end
  end
  always @(posedge clock) begin
    if(MulAddRecFNPipe_cov_write_en & MulAddRecFNPipe_cov_write_mask) begin
      MulAddRecFNPipe_cov[MulAddRecFNPipe_cov_write_addr] <= MulAddRecFNPipe_cov_write_data; // @[Coverage map for MulAddRecFNPipe]
    end
  end
endmodule
module CompareRecFN(
  input  [64:0] io_a,
  input  [64:0] io_b,
  input         io_signaling,
  output        io_lt,
  output        io_eq,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawA_sig; // @[Cat.scala 29:58]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawB_sig; // @[Cat.scala 29:58]
  wire  ordered; // @[CompareRecFN.scala 57:32]
  wire  bothInfs; // @[CompareRecFN.scala 58:33]
  wire  bothZeros; // @[CompareRecFN.scala 59:33]
  wire  eqExps; // @[CompareRecFN.scala 60:29]
  wire  _T_34; // @[CompareRecFN.scala 62:20]
  wire  _T_35; // @[CompareRecFN.scala 62:57]
  wire  _T_36; // @[CompareRecFN.scala 62:44]
  wire  common_ltMags; // @[CompareRecFN.scala 62:33]
  wire  _T_37; // @[CompareRecFN.scala 63:45]
  wire  common_eqMags; // @[CompareRecFN.scala 63:32]
  wire  _T_40; // @[CompareRecFN.scala 67:25]
  wire  _T_43; // @[CompareRecFN.scala 69:35]
  wire  _T_45; // @[CompareRecFN.scala 69:54]
  wire  _T_47; // @[CompareRecFN.scala 70:41]
  wire  _T_48; // @[CompareRecFN.scala 69:74]
  wire  _T_49; // @[CompareRecFN.scala 68:30]
  wire  _T_50; // @[CompareRecFN.scala 67:41]
  wire  ordered_lt; // @[CompareRecFN.scala 66:21]
  wire  _T_51; // @[CompareRecFN.scala 72:34]
  wire  _T_52; // @[CompareRecFN.scala 72:62]
  wire  _T_53; // @[CompareRecFN.scala 72:49]
  wire  ordered_eq; // @[CompareRecFN.scala 72:19]
  wire  _T_56; // @[common.scala 81:46]
  wire  _T_59; // @[common.scala 81:46]
  wire  _T_60; // @[CompareRecFN.scala 75:32]
  wire  _T_62; // @[CompareRecFN.scala 76:27]
  wire  invalid; // @[CompareRecFN.scala 75:58]
  wire [29:0] CompareRecFN_covSum;
  assign rawA_isZero = io_a[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_a[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_isNaN = _T_4 & io_a[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_isInf = _T_4 & ~io_a[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawA_sign = io_a[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_sExp = {1'b0,$signed(io_a[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_sig = {1'h0,~rawA_isZero,io_a[51:0]}; // @[Cat.scala 29:58]
  assign rawB_isZero = io_b[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_20 = io_b[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_isNaN = _T_20 & io_b[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_isInf = _T_20 & ~io_b[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawB_sign = io_b[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_sExp = {1'b0,$signed(io_b[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_sig = {1'h0,~rawB_isZero,io_b[51:0]}; // @[Cat.scala 29:58]
  assign ordered = ~rawA_isNaN & ~rawB_isNaN; // @[CompareRecFN.scala 57:32]
  assign bothInfs = rawA_isInf & rawB_isInf; // @[CompareRecFN.scala 58:33]
  assign bothZeros = rawA_isZero & rawB_isZero; // @[CompareRecFN.scala 59:33]
  assign eqExps = $signed(rawA_sExp) == $signed(rawB_sExp); // @[CompareRecFN.scala 60:29]
  assign _T_34 = $signed(rawA_sExp) < $signed(rawB_sExp); // @[CompareRecFN.scala 62:20]
  assign _T_35 = rawA_sig < rawB_sig; // @[CompareRecFN.scala 62:57]
  assign _T_36 = eqExps & _T_35; // @[CompareRecFN.scala 62:44]
  assign common_ltMags = _T_34 | _T_36; // @[CompareRecFN.scala 62:33]
  assign _T_37 = rawA_sig == rawB_sig; // @[CompareRecFN.scala 63:45]
  assign common_eqMags = eqExps & _T_37; // @[CompareRecFN.scala 63:32]
  assign _T_40 = rawA_sign & ~rawB_sign; // @[CompareRecFN.scala 67:25]
  assign _T_43 = rawA_sign & ~common_ltMags; // @[CompareRecFN.scala 69:35]
  assign _T_45 = _T_43 & ~common_eqMags; // @[CompareRecFN.scala 69:54]
  assign _T_47 = ~rawB_sign & common_ltMags; // @[CompareRecFN.scala 70:41]
  assign _T_48 = _T_45 | _T_47; // @[CompareRecFN.scala 69:74]
  assign _T_49 = ~bothInfs & _T_48; // @[CompareRecFN.scala 68:30]
  assign _T_50 = _T_40 | _T_49; // @[CompareRecFN.scala 67:41]
  assign ordered_lt = ~bothZeros & _T_50; // @[CompareRecFN.scala 66:21]
  assign _T_51 = rawA_sign == rawB_sign; // @[CompareRecFN.scala 72:34]
  assign _T_52 = bothInfs | common_eqMags; // @[CompareRecFN.scala 72:62]
  assign _T_53 = _T_51 & _T_52; // @[CompareRecFN.scala 72:49]
  assign ordered_eq = bothZeros | _T_53; // @[CompareRecFN.scala 72:19]
  assign _T_56 = rawA_isNaN & ~rawA_sig[51]; // @[common.scala 81:46]
  assign _T_59 = rawB_isNaN & ~rawB_sig[51]; // @[common.scala 81:46]
  assign _T_60 = _T_56 | _T_59; // @[CompareRecFN.scala 75:32]
  assign _T_62 = io_signaling & ~ordered; // @[CompareRecFN.scala 76:27]
  assign invalid = _T_60 | _T_62; // @[CompareRecFN.scala 75:58]
  assign io_lt = ordered & ordered_lt; // @[CompareRecFN.scala 78:11]
  assign io_eq = ordered & ordered_eq; // @[CompareRecFN.scala 79:11]
  assign io_exceptionFlags = {invalid,4'h0}; // @[CompareRecFN.scala 81:23]
  assign CompareRecFN_covSum = 30'h0;
  assign io_covSum = CompareRecFN_covSum;
  assign metaAssert = 1'h0;
endmodule
module RecFNToIN(
  input  [64:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_signedOut,
  output [63:0] io_out,
  output [2:0]  io_intExceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawIn_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawIn_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawIn_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawIn_sig; // @[Cat.scala 29:58]
  wire  magGeOne; // @[RecFNToIN.scala 58:30]
  wire [10:0] posExp; // @[RecFNToIN.scala 59:28]
  wire  _T_17; // @[RecFNToIN.scala 60:47]
  wire  magJustBelowOne; // @[RecFNToIN.scala 60:37]
  wire  roundingMode_near_even; // @[RecFNToIN.scala 64:53]
  wire  roundingMode_min; // @[RecFNToIN.scala 66:53]
  wire  roundingMode_max; // @[RecFNToIN.scala 67:53]
  wire  roundingMode_near_maxMag; // @[RecFNToIN.scala 68:53]
  wire  roundingMode_odd; // @[RecFNToIN.scala 69:53]
  wire [52:0] _T_19; // @[Cat.scala 29:58]
  wire [5:0] _T_21; // @[RecFNToIN.scala 81:16]
  wire [115:0] _GEN_0; // @[RecFNToIN.scala 80:50]
  wire [115:0] shiftedSig; // @[RecFNToIN.scala 80:50]
  wire  _T_24; // @[RecFNToIN.scala 86:69]
  wire [65:0] alignedSig; // @[Cat.scala 29:58]
  wire [63:0] unroundedInt; // @[RecFNToIN.scala 87:54]
  wire  _T_27; // @[RecFNToIN.scala 89:57]
  wire  common_inexact; // @[RecFNToIN.scala 89:29]
  wire  _T_30; // @[RecFNToIN.scala 91:46]
  wire  _T_32; // @[RecFNToIN.scala 91:71]
  wire  _T_33; // @[RecFNToIN.scala 91:51]
  wire  _T_34; // @[RecFNToIN.scala 91:25]
  wire  _T_37; // @[RecFNToIN.scala 92:26]
  wire  roundIncr_near_even; // @[RecFNToIN.scala 91:78]
  wire  _T_39; // @[RecFNToIN.scala 93:43]
  wire  roundIncr_near_maxMag; // @[RecFNToIN.scala 93:61]
  wire  _T_40; // @[RecFNToIN.scala 95:35]
  wire  _T_41; // @[RecFNToIN.scala 96:35]
  wire  _T_42; // @[RecFNToIN.scala 95:61]
  wire  _T_43; // @[RecFNToIN.scala 97:28]
  wire  _T_44; // @[RecFNToIN.scala 98:26]
  wire  _T_45; // @[RecFNToIN.scala 97:49]
  wire  _T_46; // @[RecFNToIN.scala 96:61]
  wire  _T_48; // @[RecFNToIN.scala 99:43]
  wire  _T_49; // @[RecFNToIN.scala 99:27]
  wire  roundIncr; // @[RecFNToIN.scala 98:46]
  wire [63:0] complUnroundedInt; // @[RecFNToIN.scala 100:32]
  wire  _T_51; // @[RecFNToIN.scala 102:23]
  wire [63:0] _T_53; // @[RecFNToIN.scala 103:31]
  wire [63:0] _T_54; // @[RecFNToIN.scala 102:12]
  wire  _T_55; // @[RecFNToIN.scala 105:31]
  wire [63:0] _GEN_1; // @[RecFNToIN.scala 105:11]
  wire [63:0] roundedInt; // @[RecFNToIN.scala 105:11]
  wire  magGeOne_atOverflowEdge; // @[RecFNToIN.scala 107:43]
  wire  _T_57; // @[RecFNToIN.scala 110:56]
  wire  roundCarryBut2; // @[RecFNToIN.scala 110:61]
  wire  _T_58; // @[RecFNToIN.scala 113:21]
  wire  _T_60; // @[RecFNToIN.scala 117:60]
  wire  _T_61; // @[RecFNToIN.scala 117:64]
  wire  _T_62; // @[RecFNToIN.scala 116:49]
  wire  _T_63; // @[RecFNToIN.scala 119:38]
  wire  _T_64; // @[RecFNToIN.scala 119:62]
  wire  _T_65; // @[RecFNToIN.scala 118:49]
  wire  _T_66; // @[RecFNToIN.scala 115:24]
  wire  _T_68; // @[RecFNToIN.scala 122:50]
  wire  _T_69; // @[RecFNToIN.scala 123:57]
  wire  _T_70; // @[RecFNToIN.scala 121:32]
  wire  _T_71; // @[RecFNToIN.scala 114:20]
  wire  _T_72; // @[RecFNToIN.scala 113:40]
  wire  _T_74; // @[RecFNToIN.scala 125:27]
  wire  _T_75; // @[RecFNToIN.scala 125:41]
  wire  common_overflow; // @[RecFNToIN.scala 112:12]
  wire  invalidExc; // @[RecFNToIN.scala 130:34]
  wire  overflow; // @[RecFNToIN.scala 131:32]
  wire  _T_79; // @[RecFNToIN.scala 132:32]
  wire  inexact; // @[RecFNToIN.scala 132:52]
  wire  excSign; // @[RecFNToIN.scala 134:32]
  wire  _T_81; // @[RecFNToIN.scala 136:27]
  wire [63:0] _T_82; // @[RecFNToIN.scala 136:12]
  wire [62:0] _T_84; // @[RecFNToIN.scala 140:12]
  wire [63:0] _GEN_2; // @[RecFNToIN.scala 139:11]
  wire [63:0] excOut; // @[RecFNToIN.scala 139:11]
  wire  _T_85; // @[RecFNToIN.scala 142:30]
  wire [1:0] _T_87; // @[Cat.scala 29:58]
  wire [29:0] RecFNToIN_covSum;
  assign rawIn_isZero = io_in[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_in[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawIn_isNaN = _T_4 & io_in[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawIn_isInf = _T_4 & ~io_in[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawIn_sign = io_in[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawIn_sExp = {1'b0,$signed(io_in[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawIn_sig = {1'h0,~rawIn_isZero,io_in[51:0]}; // @[Cat.scala 29:58]
  assign magGeOne = rawIn_sExp[11]; // @[RecFNToIN.scala 58:30]
  assign posExp = rawIn_sExp[10:0]; // @[RecFNToIN.scala 59:28]
  assign _T_17 = &posExp; // @[RecFNToIN.scala 60:47]
  assign magJustBelowOne = ~magGeOne & _T_17; // @[RecFNToIN.scala 60:37]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RecFNToIN.scala 64:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RecFNToIN.scala 66:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RecFNToIN.scala 67:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RecFNToIN.scala 68:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RecFNToIN.scala 69:53]
  assign _T_19 = {magGeOne,rawIn_sig[51:0]}; // @[Cat.scala 29:58]
  assign _T_21 = magGeOne ? rawIn_sExp[5:0] : 6'h0; // @[RecFNToIN.scala 81:16]
  assign _GEN_0 = {{63'd0}, _T_19}; // @[RecFNToIN.scala 80:50]
  assign shiftedSig = _GEN_0 << _T_21; // @[RecFNToIN.scala 80:50]
  assign _T_24 = |shiftedSig[50:0]; // @[RecFNToIN.scala 86:69]
  assign alignedSig = {shiftedSig[115:51],_T_24}; // @[Cat.scala 29:58]
  assign unroundedInt = alignedSig[65:2]; // @[RecFNToIN.scala 87:54]
  assign _T_27 = |alignedSig[1:0]; // @[RecFNToIN.scala 89:57]
  assign common_inexact = magGeOne ? _T_27 : ~rawIn_isZero; // @[RecFNToIN.scala 89:29]
  assign _T_30 = &alignedSig[2:1]; // @[RecFNToIN.scala 91:46]
  assign _T_32 = &alignedSig[1:0]; // @[RecFNToIN.scala 91:71]
  assign _T_33 = _T_30 | _T_32; // @[RecFNToIN.scala 91:51]
  assign _T_34 = magGeOne & _T_33; // @[RecFNToIN.scala 91:25]
  assign _T_37 = magJustBelowOne & _T_27; // @[RecFNToIN.scala 92:26]
  assign roundIncr_near_even = _T_34 | _T_37; // @[RecFNToIN.scala 91:78]
  assign _T_39 = magGeOne & alignedSig[1]; // @[RecFNToIN.scala 93:43]
  assign roundIncr_near_maxMag = _T_39 | magJustBelowOne; // @[RecFNToIN.scala 93:61]
  assign _T_40 = roundingMode_near_even & roundIncr_near_even; // @[RecFNToIN.scala 95:35]
  assign _T_41 = roundingMode_near_maxMag & roundIncr_near_maxMag; // @[RecFNToIN.scala 96:35]
  assign _T_42 = _T_40 | _T_41; // @[RecFNToIN.scala 95:61]
  assign _T_43 = roundingMode_min | roundingMode_odd; // @[RecFNToIN.scala 97:28]
  assign _T_44 = rawIn_sign & common_inexact; // @[RecFNToIN.scala 98:26]
  assign _T_45 = _T_43 & _T_44; // @[RecFNToIN.scala 97:49]
  assign _T_46 = _T_42 | _T_45; // @[RecFNToIN.scala 96:61]
  assign _T_48 = ~rawIn_sign & common_inexact; // @[RecFNToIN.scala 99:43]
  assign _T_49 = roundingMode_max & _T_48; // @[RecFNToIN.scala 99:27]
  assign roundIncr = _T_46 | _T_49; // @[RecFNToIN.scala 98:46]
  assign complUnroundedInt = rawIn_sign ? ~unroundedInt : unroundedInt; // @[RecFNToIN.scala 100:32]
  assign _T_51 = roundIncr ^ rawIn_sign; // @[RecFNToIN.scala 102:23]
  assign _T_53 = complUnroundedInt + 64'h1; // @[RecFNToIN.scala 103:31]
  assign _T_54 = _T_51 ? _T_53 : complUnroundedInt; // @[RecFNToIN.scala 102:12]
  assign _T_55 = roundingMode_odd & common_inexact; // @[RecFNToIN.scala 105:31]
  assign _GEN_1 = {{63'd0}, _T_55}; // @[RecFNToIN.scala 105:11]
  assign roundedInt = _T_54 | _GEN_1; // @[RecFNToIN.scala 105:11]
  assign magGeOne_atOverflowEdge = posExp == 11'h3f; // @[RecFNToIN.scala 107:43]
  assign _T_57 = &unroundedInt[61:0]; // @[RecFNToIN.scala 110:56]
  assign roundCarryBut2 = _T_57 & roundIncr; // @[RecFNToIN.scala 110:61]
  assign _T_58 = posExp >= 11'h40; // @[RecFNToIN.scala 113:21]
  assign _T_60 = |unroundedInt[62:0]; // @[RecFNToIN.scala 117:60]
  assign _T_61 = _T_60 | roundIncr; // @[RecFNToIN.scala 117:64]
  assign _T_62 = magGeOne_atOverflowEdge & _T_61; // @[RecFNToIN.scala 116:49]
  assign _T_63 = posExp == 11'h3e; // @[RecFNToIN.scala 119:38]
  assign _T_64 = _T_63 & roundCarryBut2; // @[RecFNToIN.scala 119:62]
  assign _T_65 = magGeOne_atOverflowEdge | _T_64; // @[RecFNToIN.scala 118:49]
  assign _T_66 = rawIn_sign ? _T_62 : _T_65; // @[RecFNToIN.scala 115:24]
  assign _T_68 = magGeOne_atOverflowEdge & unroundedInt[62]; // @[RecFNToIN.scala 122:50]
  assign _T_69 = _T_68 & roundCarryBut2; // @[RecFNToIN.scala 123:57]
  assign _T_70 = rawIn_sign | _T_69; // @[RecFNToIN.scala 121:32]
  assign _T_71 = io_signedOut ? _T_66 : _T_70; // @[RecFNToIN.scala 114:20]
  assign _T_72 = _T_58 | _T_71; // @[RecFNToIN.scala 113:40]
  assign _T_74 = ~io_signedOut & rawIn_sign; // @[RecFNToIN.scala 125:27]
  assign _T_75 = _T_74 & roundIncr; // @[RecFNToIN.scala 125:41]
  assign common_overflow = magGeOne ? _T_72 : _T_75; // @[RecFNToIN.scala 112:12]
  assign invalidExc = rawIn_isNaN | rawIn_isInf; // @[RecFNToIN.scala 130:34]
  assign overflow = ~invalidExc & common_overflow; // @[RecFNToIN.scala 131:32]
  assign _T_79 = ~invalidExc & ~common_overflow; // @[RecFNToIN.scala 132:32]
  assign inexact = _T_79 & common_inexact; // @[RecFNToIN.scala 132:52]
  assign excSign = ~rawIn_isNaN & rawIn_sign; // @[RecFNToIN.scala 134:32]
  assign _T_81 = io_signedOut == excSign; // @[RecFNToIN.scala 136:27]
  assign _T_82 = _T_81 ? 64'h8000000000000000 : 64'h0; // @[RecFNToIN.scala 136:12]
  assign _T_84 = excSign ? 63'h0 : 63'h7fffffffffffffff; // @[RecFNToIN.scala 140:12]
  assign _GEN_2 = {{1'd0}, _T_84}; // @[RecFNToIN.scala 139:11]
  assign excOut = _T_82 | _GEN_2; // @[RecFNToIN.scala 139:11]
  assign _T_85 = invalidExc | common_overflow; // @[RecFNToIN.scala 142:30]
  assign _T_87 = {invalidExc,overflow}; // @[Cat.scala 29:58]
  assign io_out = _T_85 ? excOut : roundedInt; // @[RecFNToIN.scala 142:12]
  assign io_intExceptionFlags = {_T_87,inexact}; // @[RecFNToIN.scala 143:26]
  assign RecFNToIN_covSum = 30'h0;
  assign io_covSum = RecFNToIN_covSum;
  assign metaAssert = 1'h0;
endmodule
module RecFNToIN_1(
  input  [64:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_signedOut,
  output [2:0]  io_intExceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawIn_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawIn_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawIn_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawIn_sig; // @[Cat.scala 29:58]
  wire  magGeOne; // @[RecFNToIN.scala 58:30]
  wire [10:0] posExp; // @[RecFNToIN.scala 59:28]
  wire  _T_17; // @[RecFNToIN.scala 60:47]
  wire  magJustBelowOne; // @[RecFNToIN.scala 60:37]
  wire  roundingMode_near_even; // @[RecFNToIN.scala 64:53]
  wire  roundingMode_min; // @[RecFNToIN.scala 66:53]
  wire  roundingMode_max; // @[RecFNToIN.scala 67:53]
  wire  roundingMode_near_maxMag; // @[RecFNToIN.scala 68:53]
  wire  roundingMode_odd; // @[RecFNToIN.scala 69:53]
  wire [52:0] _T_19; // @[Cat.scala 29:58]
  wire [4:0] _T_21; // @[RecFNToIN.scala 81:16]
  wire [83:0] _GEN_0; // @[RecFNToIN.scala 80:50]
  wire [83:0] shiftedSig; // @[RecFNToIN.scala 80:50]
  wire  _T_24; // @[RecFNToIN.scala 86:69]
  wire [33:0] alignedSig; // @[Cat.scala 29:58]
  wire [31:0] unroundedInt; // @[RecFNToIN.scala 87:54]
  wire  _T_27; // @[RecFNToIN.scala 89:57]
  wire  common_inexact; // @[RecFNToIN.scala 89:29]
  wire  _T_30; // @[RecFNToIN.scala 91:46]
  wire  _T_32; // @[RecFNToIN.scala 91:71]
  wire  _T_33; // @[RecFNToIN.scala 91:51]
  wire  _T_34; // @[RecFNToIN.scala 91:25]
  wire  _T_37; // @[RecFNToIN.scala 92:26]
  wire  roundIncr_near_even; // @[RecFNToIN.scala 91:78]
  wire  _T_39; // @[RecFNToIN.scala 93:43]
  wire  roundIncr_near_maxMag; // @[RecFNToIN.scala 93:61]
  wire  _T_40; // @[RecFNToIN.scala 95:35]
  wire  _T_41; // @[RecFNToIN.scala 96:35]
  wire  _T_42; // @[RecFNToIN.scala 95:61]
  wire  _T_43; // @[RecFNToIN.scala 97:28]
  wire  _T_44; // @[RecFNToIN.scala 98:26]
  wire  _T_45; // @[RecFNToIN.scala 97:49]
  wire  _T_46; // @[RecFNToIN.scala 96:61]
  wire  _T_48; // @[RecFNToIN.scala 99:43]
  wire  _T_49; // @[RecFNToIN.scala 99:27]
  wire  roundIncr; // @[RecFNToIN.scala 98:46]
  wire  magGeOne_atOverflowEdge; // @[RecFNToIN.scala 107:43]
  wire  _T_57; // @[RecFNToIN.scala 110:56]
  wire  roundCarryBut2; // @[RecFNToIN.scala 110:61]
  wire  _T_58; // @[RecFNToIN.scala 113:21]
  wire  _T_60; // @[RecFNToIN.scala 117:60]
  wire  _T_61; // @[RecFNToIN.scala 117:64]
  wire  _T_62; // @[RecFNToIN.scala 116:49]
  wire  _T_63; // @[RecFNToIN.scala 119:38]
  wire  _T_64; // @[RecFNToIN.scala 119:62]
  wire  _T_65; // @[RecFNToIN.scala 118:49]
  wire  _T_66; // @[RecFNToIN.scala 115:24]
  wire  _T_68; // @[RecFNToIN.scala 122:50]
  wire  _T_69; // @[RecFNToIN.scala 123:57]
  wire  _T_70; // @[RecFNToIN.scala 121:32]
  wire  _T_71; // @[RecFNToIN.scala 114:20]
  wire  _T_72; // @[RecFNToIN.scala 113:40]
  wire  _T_74; // @[RecFNToIN.scala 125:27]
  wire  _T_75; // @[RecFNToIN.scala 125:41]
  wire  common_overflow; // @[RecFNToIN.scala 112:12]
  wire  invalidExc; // @[RecFNToIN.scala 130:34]
  wire  overflow; // @[RecFNToIN.scala 131:32]
  wire  _T_79; // @[RecFNToIN.scala 132:32]
  wire  inexact; // @[RecFNToIN.scala 132:52]
  wire [1:0] _T_87; // @[Cat.scala 29:58]
  wire [29:0] RecFNToIN_1_covSum;
  assign rawIn_isZero = io_in[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_in[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawIn_isNaN = _T_4 & io_in[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawIn_isInf = _T_4 & ~io_in[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawIn_sign = io_in[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawIn_sExp = {1'b0,$signed(io_in[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawIn_sig = {1'h0,~rawIn_isZero,io_in[51:0]}; // @[Cat.scala 29:58]
  assign magGeOne = rawIn_sExp[11]; // @[RecFNToIN.scala 58:30]
  assign posExp = rawIn_sExp[10:0]; // @[RecFNToIN.scala 59:28]
  assign _T_17 = &posExp; // @[RecFNToIN.scala 60:47]
  assign magJustBelowOne = ~magGeOne & _T_17; // @[RecFNToIN.scala 60:37]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RecFNToIN.scala 64:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RecFNToIN.scala 66:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RecFNToIN.scala 67:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RecFNToIN.scala 68:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RecFNToIN.scala 69:53]
  assign _T_19 = {magGeOne,rawIn_sig[51:0]}; // @[Cat.scala 29:58]
  assign _T_21 = magGeOne ? rawIn_sExp[4:0] : 5'h0; // @[RecFNToIN.scala 81:16]
  assign _GEN_0 = {{31'd0}, _T_19}; // @[RecFNToIN.scala 80:50]
  assign shiftedSig = _GEN_0 << _T_21; // @[RecFNToIN.scala 80:50]
  assign _T_24 = |shiftedSig[50:0]; // @[RecFNToIN.scala 86:69]
  assign alignedSig = {shiftedSig[83:51],_T_24}; // @[Cat.scala 29:58]
  assign unroundedInt = alignedSig[33:2]; // @[RecFNToIN.scala 87:54]
  assign _T_27 = |alignedSig[1:0]; // @[RecFNToIN.scala 89:57]
  assign common_inexact = magGeOne ? _T_27 : ~rawIn_isZero; // @[RecFNToIN.scala 89:29]
  assign _T_30 = &alignedSig[2:1]; // @[RecFNToIN.scala 91:46]
  assign _T_32 = &alignedSig[1:0]; // @[RecFNToIN.scala 91:71]
  assign _T_33 = _T_30 | _T_32; // @[RecFNToIN.scala 91:51]
  assign _T_34 = magGeOne & _T_33; // @[RecFNToIN.scala 91:25]
  assign _T_37 = magJustBelowOne & _T_27; // @[RecFNToIN.scala 92:26]
  assign roundIncr_near_even = _T_34 | _T_37; // @[RecFNToIN.scala 91:78]
  assign _T_39 = magGeOne & alignedSig[1]; // @[RecFNToIN.scala 93:43]
  assign roundIncr_near_maxMag = _T_39 | magJustBelowOne; // @[RecFNToIN.scala 93:61]
  assign _T_40 = roundingMode_near_even & roundIncr_near_even; // @[RecFNToIN.scala 95:35]
  assign _T_41 = roundingMode_near_maxMag & roundIncr_near_maxMag; // @[RecFNToIN.scala 96:35]
  assign _T_42 = _T_40 | _T_41; // @[RecFNToIN.scala 95:61]
  assign _T_43 = roundingMode_min | roundingMode_odd; // @[RecFNToIN.scala 97:28]
  assign _T_44 = rawIn_sign & common_inexact; // @[RecFNToIN.scala 98:26]
  assign _T_45 = _T_43 & _T_44; // @[RecFNToIN.scala 97:49]
  assign _T_46 = _T_42 | _T_45; // @[RecFNToIN.scala 96:61]
  assign _T_48 = ~rawIn_sign & common_inexact; // @[RecFNToIN.scala 99:43]
  assign _T_49 = roundingMode_max & _T_48; // @[RecFNToIN.scala 99:27]
  assign roundIncr = _T_46 | _T_49; // @[RecFNToIN.scala 98:46]
  assign magGeOne_atOverflowEdge = posExp == 11'h1f; // @[RecFNToIN.scala 107:43]
  assign _T_57 = &unroundedInt[29:0]; // @[RecFNToIN.scala 110:56]
  assign roundCarryBut2 = _T_57 & roundIncr; // @[RecFNToIN.scala 110:61]
  assign _T_58 = posExp >= 11'h20; // @[RecFNToIN.scala 113:21]
  assign _T_60 = |unroundedInt[30:0]; // @[RecFNToIN.scala 117:60]
  assign _T_61 = _T_60 | roundIncr; // @[RecFNToIN.scala 117:64]
  assign _T_62 = magGeOne_atOverflowEdge & _T_61; // @[RecFNToIN.scala 116:49]
  assign _T_63 = posExp == 11'h1e; // @[RecFNToIN.scala 119:38]
  assign _T_64 = _T_63 & roundCarryBut2; // @[RecFNToIN.scala 119:62]
  assign _T_65 = magGeOne_atOverflowEdge | _T_64; // @[RecFNToIN.scala 118:49]
  assign _T_66 = rawIn_sign ? _T_62 : _T_65; // @[RecFNToIN.scala 115:24]
  assign _T_68 = magGeOne_atOverflowEdge & unroundedInt[30]; // @[RecFNToIN.scala 122:50]
  assign _T_69 = _T_68 & roundCarryBut2; // @[RecFNToIN.scala 123:57]
  assign _T_70 = rawIn_sign | _T_69; // @[RecFNToIN.scala 121:32]
  assign _T_71 = io_signedOut ? _T_66 : _T_70; // @[RecFNToIN.scala 114:20]
  assign _T_72 = _T_58 | _T_71; // @[RecFNToIN.scala 113:40]
  assign _T_74 = ~io_signedOut & rawIn_sign; // @[RecFNToIN.scala 125:27]
  assign _T_75 = _T_74 & roundIncr; // @[RecFNToIN.scala 125:41]
  assign common_overflow = magGeOne ? _T_72 : _T_75; // @[RecFNToIN.scala 112:12]
  assign invalidExc = rawIn_isNaN | rawIn_isInf; // @[RecFNToIN.scala 130:34]
  assign overflow = ~invalidExc & common_overflow; // @[RecFNToIN.scala 131:32]
  assign _T_79 = ~invalidExc & ~common_overflow; // @[RecFNToIN.scala 132:32]
  assign inexact = _T_79 & common_inexact; // @[RecFNToIN.scala 132:52]
  assign _T_87 = {invalidExc,overflow}; // @[Cat.scala 29:58]
  assign io_intExceptionFlags = {_T_87,inexact}; // @[RecFNToIN.scala 143:26]
  assign RecFNToIN_1_covSum = 30'h0;
  assign io_covSum = RecFNToIN_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module INToRecFN(
  input         io_signedIn,
  input  [63:0] io_in,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[INToRecFN.scala 59:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[INToRecFN.scala 59:15]
  wire [8:0] roundAnyRawFNToRecFN_io_in_sExp; // @[INToRecFN.scala 59:15]
  wire [64:0] roundAnyRawFNToRecFN_io_in_sig; // @[INToRecFN.scala 59:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[INToRecFN.scala 59:15]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 59:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 59:15]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[INToRecFN.scala 59:15]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[INToRecFN.scala 59:15]
  wire  intAsRawFloat_sign; // @[rawFloatFromIN.scala 50:29]
  wire [63:0] _T_3; // @[rawFloatFromIN.scala 51:31]
  wire [63:0] _T_4; // @[rawFloatFromIN.scala 51:24]
  wire [127:0] _T_5; // @[Cat.scala 29:58]
  wire [5:0] _T_71; // @[Mux.scala 47:69]
  wire [5:0] _T_72; // @[Mux.scala 47:69]
  wire [5:0] _T_73; // @[Mux.scala 47:69]
  wire [5:0] _T_74; // @[Mux.scala 47:69]
  wire [5:0] _T_75; // @[Mux.scala 47:69]
  wire [5:0] _T_76; // @[Mux.scala 47:69]
  wire [5:0] _T_77; // @[Mux.scala 47:69]
  wire [5:0] _T_78; // @[Mux.scala 47:69]
  wire [5:0] _T_79; // @[Mux.scala 47:69]
  wire [5:0] _T_80; // @[Mux.scala 47:69]
  wire [5:0] _T_81; // @[Mux.scala 47:69]
  wire [5:0] _T_82; // @[Mux.scala 47:69]
  wire [5:0] _T_83; // @[Mux.scala 47:69]
  wire [5:0] _T_84; // @[Mux.scala 47:69]
  wire [5:0] _T_85; // @[Mux.scala 47:69]
  wire [5:0] _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_106; // @[Mux.scala 47:69]
  wire [5:0] _T_107; // @[Mux.scala 47:69]
  wire [5:0] _T_108; // @[Mux.scala 47:69]
  wire [5:0] _T_109; // @[Mux.scala 47:69]
  wire [5:0] _T_110; // @[Mux.scala 47:69]
  wire [5:0] _T_111; // @[Mux.scala 47:69]
  wire [5:0] _T_112; // @[Mux.scala 47:69]
  wire [5:0] _T_113; // @[Mux.scala 47:69]
  wire [5:0] _T_114; // @[Mux.scala 47:69]
  wire [5:0] _T_115; // @[Mux.scala 47:69]
  wire [5:0] _T_116; // @[Mux.scala 47:69]
  wire [5:0] _T_117; // @[Mux.scala 47:69]
  wire [5:0] _T_118; // @[Mux.scala 47:69]
  wire [5:0] _T_119; // @[Mux.scala 47:69]
  wire [5:0] _T_120; // @[Mux.scala 47:69]
  wire [5:0] _T_121; // @[Mux.scala 47:69]
  wire [5:0] _T_122; // @[Mux.scala 47:69]
  wire [5:0] _T_123; // @[Mux.scala 47:69]
  wire [5:0] _T_124; // @[Mux.scala 47:69]
  wire [5:0] _T_125; // @[Mux.scala 47:69]
  wire [5:0] _T_126; // @[Mux.scala 47:69]
  wire [5:0] _T_127; // @[Mux.scala 47:69]
  wire [5:0] _T_128; // @[Mux.scala 47:69]
  wire [5:0] _T_129; // @[Mux.scala 47:69]
  wire [5:0] _T_130; // @[Mux.scala 47:69]
  wire [5:0] _T_131; // @[Mux.scala 47:69]
  wire [5:0] _T_132; // @[Mux.scala 47:69]
  wire [5:0] _T_133; // @[Mux.scala 47:69]
  wire [126:0] _GEN_0; // @[rawFloatFromIN.scala 55:22]
  wire [126:0] _T_134; // @[rawFloatFromIN.scala 55:22]
  wire [7:0] _T_140; // @[Cat.scala 29:58]
  wire [29:0] INToRecFN_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_1 roundAnyRawFNToRecFN ( // @[INToRecFN.scala 59:15]
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign intAsRawFloat_sign = io_signedIn & io_in[63]; // @[rawFloatFromIN.scala 50:29]
  assign _T_3 = 64'h0 - io_in; // @[rawFloatFromIN.scala 51:31]
  assign _T_4 = intAsRawFloat_sign ? _T_3 : io_in; // @[rawFloatFromIN.scala 51:24]
  assign _T_5 = {64'h0,_T_4}; // @[Cat.scala 29:58]
  assign _T_71 = _T_5[1] ? 6'h3e : 6'h3f; // @[Mux.scala 47:69]
  assign _T_72 = _T_5[2] ? 6'h3d : _T_71; // @[Mux.scala 47:69]
  assign _T_73 = _T_5[3] ? 6'h3c : _T_72; // @[Mux.scala 47:69]
  assign _T_74 = _T_5[4] ? 6'h3b : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = _T_5[5] ? 6'h3a : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = _T_5[6] ? 6'h39 : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = _T_5[7] ? 6'h38 : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = _T_5[8] ? 6'h37 : _T_77; // @[Mux.scala 47:69]
  assign _T_79 = _T_5[9] ? 6'h36 : _T_78; // @[Mux.scala 47:69]
  assign _T_80 = _T_5[10] ? 6'h35 : _T_79; // @[Mux.scala 47:69]
  assign _T_81 = _T_5[11] ? 6'h34 : _T_80; // @[Mux.scala 47:69]
  assign _T_82 = _T_5[12] ? 6'h33 : _T_81; // @[Mux.scala 47:69]
  assign _T_83 = _T_5[13] ? 6'h32 : _T_82; // @[Mux.scala 47:69]
  assign _T_84 = _T_5[14] ? 6'h31 : _T_83; // @[Mux.scala 47:69]
  assign _T_85 = _T_5[15] ? 6'h30 : _T_84; // @[Mux.scala 47:69]
  assign _T_86 = _T_5[16] ? 6'h2f : _T_85; // @[Mux.scala 47:69]
  assign _T_87 = _T_5[17] ? 6'h2e : _T_86; // @[Mux.scala 47:69]
  assign _T_88 = _T_5[18] ? 6'h2d : _T_87; // @[Mux.scala 47:69]
  assign _T_89 = _T_5[19] ? 6'h2c : _T_88; // @[Mux.scala 47:69]
  assign _T_90 = _T_5[20] ? 6'h2b : _T_89; // @[Mux.scala 47:69]
  assign _T_91 = _T_5[21] ? 6'h2a : _T_90; // @[Mux.scala 47:69]
  assign _T_92 = _T_5[22] ? 6'h29 : _T_91; // @[Mux.scala 47:69]
  assign _T_93 = _T_5[23] ? 6'h28 : _T_92; // @[Mux.scala 47:69]
  assign _T_94 = _T_5[24] ? 6'h27 : _T_93; // @[Mux.scala 47:69]
  assign _T_95 = _T_5[25] ? 6'h26 : _T_94; // @[Mux.scala 47:69]
  assign _T_96 = _T_5[26] ? 6'h25 : _T_95; // @[Mux.scala 47:69]
  assign _T_97 = _T_5[27] ? 6'h24 : _T_96; // @[Mux.scala 47:69]
  assign _T_98 = _T_5[28] ? 6'h23 : _T_97; // @[Mux.scala 47:69]
  assign _T_99 = _T_5[29] ? 6'h22 : _T_98; // @[Mux.scala 47:69]
  assign _T_100 = _T_5[30] ? 6'h21 : _T_99; // @[Mux.scala 47:69]
  assign _T_101 = _T_5[31] ? 6'h20 : _T_100; // @[Mux.scala 47:69]
  assign _T_102 = _T_5[32] ? 6'h1f : _T_101; // @[Mux.scala 47:69]
  assign _T_103 = _T_5[33] ? 6'h1e : _T_102; // @[Mux.scala 47:69]
  assign _T_104 = _T_5[34] ? 6'h1d : _T_103; // @[Mux.scala 47:69]
  assign _T_105 = _T_5[35] ? 6'h1c : _T_104; // @[Mux.scala 47:69]
  assign _T_106 = _T_5[36] ? 6'h1b : _T_105; // @[Mux.scala 47:69]
  assign _T_107 = _T_5[37] ? 6'h1a : _T_106; // @[Mux.scala 47:69]
  assign _T_108 = _T_5[38] ? 6'h19 : _T_107; // @[Mux.scala 47:69]
  assign _T_109 = _T_5[39] ? 6'h18 : _T_108; // @[Mux.scala 47:69]
  assign _T_110 = _T_5[40] ? 6'h17 : _T_109; // @[Mux.scala 47:69]
  assign _T_111 = _T_5[41] ? 6'h16 : _T_110; // @[Mux.scala 47:69]
  assign _T_112 = _T_5[42] ? 6'h15 : _T_111; // @[Mux.scala 47:69]
  assign _T_113 = _T_5[43] ? 6'h14 : _T_112; // @[Mux.scala 47:69]
  assign _T_114 = _T_5[44] ? 6'h13 : _T_113; // @[Mux.scala 47:69]
  assign _T_115 = _T_5[45] ? 6'h12 : _T_114; // @[Mux.scala 47:69]
  assign _T_116 = _T_5[46] ? 6'h11 : _T_115; // @[Mux.scala 47:69]
  assign _T_117 = _T_5[47] ? 6'h10 : _T_116; // @[Mux.scala 47:69]
  assign _T_118 = _T_5[48] ? 6'hf : _T_117; // @[Mux.scala 47:69]
  assign _T_119 = _T_5[49] ? 6'he : _T_118; // @[Mux.scala 47:69]
  assign _T_120 = _T_5[50] ? 6'hd : _T_119; // @[Mux.scala 47:69]
  assign _T_121 = _T_5[51] ? 6'hc : _T_120; // @[Mux.scala 47:69]
  assign _T_122 = _T_5[52] ? 6'hb : _T_121; // @[Mux.scala 47:69]
  assign _T_123 = _T_5[53] ? 6'ha : _T_122; // @[Mux.scala 47:69]
  assign _T_124 = _T_5[54] ? 6'h9 : _T_123; // @[Mux.scala 47:69]
  assign _T_125 = _T_5[55] ? 6'h8 : _T_124; // @[Mux.scala 47:69]
  assign _T_126 = _T_5[56] ? 6'h7 : _T_125; // @[Mux.scala 47:69]
  assign _T_127 = _T_5[57] ? 6'h6 : _T_126; // @[Mux.scala 47:69]
  assign _T_128 = _T_5[58] ? 6'h5 : _T_127; // @[Mux.scala 47:69]
  assign _T_129 = _T_5[59] ? 6'h4 : _T_128; // @[Mux.scala 47:69]
  assign _T_130 = _T_5[60] ? 6'h3 : _T_129; // @[Mux.scala 47:69]
  assign _T_131 = _T_5[61] ? 6'h2 : _T_130; // @[Mux.scala 47:69]
  assign _T_132 = _T_5[62] ? 6'h1 : _T_131; // @[Mux.scala 47:69]
  assign _T_133 = _T_5[63] ? 6'h0 : _T_132; // @[Mux.scala 47:69]
  assign _GEN_0 = {{63'd0}, _T_5[63:0]}; // @[rawFloatFromIN.scala 55:22]
  assign _T_134 = _GEN_0 << _T_133; // @[rawFloatFromIN.scala 55:22]
  assign _T_140 = {2'h2,~_T_133}; // @[Cat.scala 29:58]
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 72:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 73:23]
  assign roundAnyRawFNToRecFN_io_in_isZero = ~_T_134[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_signedIn & io_in[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(_T_140)}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sig = {{1'd0}, _T_134[63:0]}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[INToRecFN.scala 70:44]
  assign INToRecFN_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = INToRecFN_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module INToRecFN_1(
  input         io_signedIn,
  input  [63:0] io_in,
  input  [2:0]  io_roundingMode,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[INToRecFN.scala 59:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[INToRecFN.scala 59:15]
  wire [8:0] roundAnyRawFNToRecFN_io_in_sExp; // @[INToRecFN.scala 59:15]
  wire [64:0] roundAnyRawFNToRecFN_io_in_sig; // @[INToRecFN.scala 59:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[INToRecFN.scala 59:15]
  wire [64:0] roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 59:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 59:15]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[INToRecFN.scala 59:15]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[INToRecFN.scala 59:15]
  wire  intAsRawFloat_sign; // @[rawFloatFromIN.scala 50:29]
  wire [63:0] _T_3; // @[rawFloatFromIN.scala 51:31]
  wire [63:0] _T_4; // @[rawFloatFromIN.scala 51:24]
  wire [127:0] _T_5; // @[Cat.scala 29:58]
  wire [5:0] _T_71; // @[Mux.scala 47:69]
  wire [5:0] _T_72; // @[Mux.scala 47:69]
  wire [5:0] _T_73; // @[Mux.scala 47:69]
  wire [5:0] _T_74; // @[Mux.scala 47:69]
  wire [5:0] _T_75; // @[Mux.scala 47:69]
  wire [5:0] _T_76; // @[Mux.scala 47:69]
  wire [5:0] _T_77; // @[Mux.scala 47:69]
  wire [5:0] _T_78; // @[Mux.scala 47:69]
  wire [5:0] _T_79; // @[Mux.scala 47:69]
  wire [5:0] _T_80; // @[Mux.scala 47:69]
  wire [5:0] _T_81; // @[Mux.scala 47:69]
  wire [5:0] _T_82; // @[Mux.scala 47:69]
  wire [5:0] _T_83; // @[Mux.scala 47:69]
  wire [5:0] _T_84; // @[Mux.scala 47:69]
  wire [5:0] _T_85; // @[Mux.scala 47:69]
  wire [5:0] _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_106; // @[Mux.scala 47:69]
  wire [5:0] _T_107; // @[Mux.scala 47:69]
  wire [5:0] _T_108; // @[Mux.scala 47:69]
  wire [5:0] _T_109; // @[Mux.scala 47:69]
  wire [5:0] _T_110; // @[Mux.scala 47:69]
  wire [5:0] _T_111; // @[Mux.scala 47:69]
  wire [5:0] _T_112; // @[Mux.scala 47:69]
  wire [5:0] _T_113; // @[Mux.scala 47:69]
  wire [5:0] _T_114; // @[Mux.scala 47:69]
  wire [5:0] _T_115; // @[Mux.scala 47:69]
  wire [5:0] _T_116; // @[Mux.scala 47:69]
  wire [5:0] _T_117; // @[Mux.scala 47:69]
  wire [5:0] _T_118; // @[Mux.scala 47:69]
  wire [5:0] _T_119; // @[Mux.scala 47:69]
  wire [5:0] _T_120; // @[Mux.scala 47:69]
  wire [5:0] _T_121; // @[Mux.scala 47:69]
  wire [5:0] _T_122; // @[Mux.scala 47:69]
  wire [5:0] _T_123; // @[Mux.scala 47:69]
  wire [5:0] _T_124; // @[Mux.scala 47:69]
  wire [5:0] _T_125; // @[Mux.scala 47:69]
  wire [5:0] _T_126; // @[Mux.scala 47:69]
  wire [5:0] _T_127; // @[Mux.scala 47:69]
  wire [5:0] _T_128; // @[Mux.scala 47:69]
  wire [5:0] _T_129; // @[Mux.scala 47:69]
  wire [5:0] _T_130; // @[Mux.scala 47:69]
  wire [5:0] _T_131; // @[Mux.scala 47:69]
  wire [5:0] _T_132; // @[Mux.scala 47:69]
  wire [5:0] _T_133; // @[Mux.scala 47:69]
  wire [126:0] _GEN_0; // @[rawFloatFromIN.scala 55:22]
  wire [126:0] _T_134; // @[rawFloatFromIN.scala 55:22]
  wire [7:0] _T_140; // @[Cat.scala 29:58]
  wire [29:0] INToRecFN_1_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_2 roundAnyRawFNToRecFN ( // @[INToRecFN.scala 59:15]
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign intAsRawFloat_sign = io_signedIn & io_in[63]; // @[rawFloatFromIN.scala 50:29]
  assign _T_3 = 64'h0 - io_in; // @[rawFloatFromIN.scala 51:31]
  assign _T_4 = intAsRawFloat_sign ? _T_3 : io_in; // @[rawFloatFromIN.scala 51:24]
  assign _T_5 = {64'h0,_T_4}; // @[Cat.scala 29:58]
  assign _T_71 = _T_5[1] ? 6'h3e : 6'h3f; // @[Mux.scala 47:69]
  assign _T_72 = _T_5[2] ? 6'h3d : _T_71; // @[Mux.scala 47:69]
  assign _T_73 = _T_5[3] ? 6'h3c : _T_72; // @[Mux.scala 47:69]
  assign _T_74 = _T_5[4] ? 6'h3b : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = _T_5[5] ? 6'h3a : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = _T_5[6] ? 6'h39 : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = _T_5[7] ? 6'h38 : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = _T_5[8] ? 6'h37 : _T_77; // @[Mux.scala 47:69]
  assign _T_79 = _T_5[9] ? 6'h36 : _T_78; // @[Mux.scala 47:69]
  assign _T_80 = _T_5[10] ? 6'h35 : _T_79; // @[Mux.scala 47:69]
  assign _T_81 = _T_5[11] ? 6'h34 : _T_80; // @[Mux.scala 47:69]
  assign _T_82 = _T_5[12] ? 6'h33 : _T_81; // @[Mux.scala 47:69]
  assign _T_83 = _T_5[13] ? 6'h32 : _T_82; // @[Mux.scala 47:69]
  assign _T_84 = _T_5[14] ? 6'h31 : _T_83; // @[Mux.scala 47:69]
  assign _T_85 = _T_5[15] ? 6'h30 : _T_84; // @[Mux.scala 47:69]
  assign _T_86 = _T_5[16] ? 6'h2f : _T_85; // @[Mux.scala 47:69]
  assign _T_87 = _T_5[17] ? 6'h2e : _T_86; // @[Mux.scala 47:69]
  assign _T_88 = _T_5[18] ? 6'h2d : _T_87; // @[Mux.scala 47:69]
  assign _T_89 = _T_5[19] ? 6'h2c : _T_88; // @[Mux.scala 47:69]
  assign _T_90 = _T_5[20] ? 6'h2b : _T_89; // @[Mux.scala 47:69]
  assign _T_91 = _T_5[21] ? 6'h2a : _T_90; // @[Mux.scala 47:69]
  assign _T_92 = _T_5[22] ? 6'h29 : _T_91; // @[Mux.scala 47:69]
  assign _T_93 = _T_5[23] ? 6'h28 : _T_92; // @[Mux.scala 47:69]
  assign _T_94 = _T_5[24] ? 6'h27 : _T_93; // @[Mux.scala 47:69]
  assign _T_95 = _T_5[25] ? 6'h26 : _T_94; // @[Mux.scala 47:69]
  assign _T_96 = _T_5[26] ? 6'h25 : _T_95; // @[Mux.scala 47:69]
  assign _T_97 = _T_5[27] ? 6'h24 : _T_96; // @[Mux.scala 47:69]
  assign _T_98 = _T_5[28] ? 6'h23 : _T_97; // @[Mux.scala 47:69]
  assign _T_99 = _T_5[29] ? 6'h22 : _T_98; // @[Mux.scala 47:69]
  assign _T_100 = _T_5[30] ? 6'h21 : _T_99; // @[Mux.scala 47:69]
  assign _T_101 = _T_5[31] ? 6'h20 : _T_100; // @[Mux.scala 47:69]
  assign _T_102 = _T_5[32] ? 6'h1f : _T_101; // @[Mux.scala 47:69]
  assign _T_103 = _T_5[33] ? 6'h1e : _T_102; // @[Mux.scala 47:69]
  assign _T_104 = _T_5[34] ? 6'h1d : _T_103; // @[Mux.scala 47:69]
  assign _T_105 = _T_5[35] ? 6'h1c : _T_104; // @[Mux.scala 47:69]
  assign _T_106 = _T_5[36] ? 6'h1b : _T_105; // @[Mux.scala 47:69]
  assign _T_107 = _T_5[37] ? 6'h1a : _T_106; // @[Mux.scala 47:69]
  assign _T_108 = _T_5[38] ? 6'h19 : _T_107; // @[Mux.scala 47:69]
  assign _T_109 = _T_5[39] ? 6'h18 : _T_108; // @[Mux.scala 47:69]
  assign _T_110 = _T_5[40] ? 6'h17 : _T_109; // @[Mux.scala 47:69]
  assign _T_111 = _T_5[41] ? 6'h16 : _T_110; // @[Mux.scala 47:69]
  assign _T_112 = _T_5[42] ? 6'h15 : _T_111; // @[Mux.scala 47:69]
  assign _T_113 = _T_5[43] ? 6'h14 : _T_112; // @[Mux.scala 47:69]
  assign _T_114 = _T_5[44] ? 6'h13 : _T_113; // @[Mux.scala 47:69]
  assign _T_115 = _T_5[45] ? 6'h12 : _T_114; // @[Mux.scala 47:69]
  assign _T_116 = _T_5[46] ? 6'h11 : _T_115; // @[Mux.scala 47:69]
  assign _T_117 = _T_5[47] ? 6'h10 : _T_116; // @[Mux.scala 47:69]
  assign _T_118 = _T_5[48] ? 6'hf : _T_117; // @[Mux.scala 47:69]
  assign _T_119 = _T_5[49] ? 6'he : _T_118; // @[Mux.scala 47:69]
  assign _T_120 = _T_5[50] ? 6'hd : _T_119; // @[Mux.scala 47:69]
  assign _T_121 = _T_5[51] ? 6'hc : _T_120; // @[Mux.scala 47:69]
  assign _T_122 = _T_5[52] ? 6'hb : _T_121; // @[Mux.scala 47:69]
  assign _T_123 = _T_5[53] ? 6'ha : _T_122; // @[Mux.scala 47:69]
  assign _T_124 = _T_5[54] ? 6'h9 : _T_123; // @[Mux.scala 47:69]
  assign _T_125 = _T_5[55] ? 6'h8 : _T_124; // @[Mux.scala 47:69]
  assign _T_126 = _T_5[56] ? 6'h7 : _T_125; // @[Mux.scala 47:69]
  assign _T_127 = _T_5[57] ? 6'h6 : _T_126; // @[Mux.scala 47:69]
  assign _T_128 = _T_5[58] ? 6'h5 : _T_127; // @[Mux.scala 47:69]
  assign _T_129 = _T_5[59] ? 6'h4 : _T_128; // @[Mux.scala 47:69]
  assign _T_130 = _T_5[60] ? 6'h3 : _T_129; // @[Mux.scala 47:69]
  assign _T_131 = _T_5[61] ? 6'h2 : _T_130; // @[Mux.scala 47:69]
  assign _T_132 = _T_5[62] ? 6'h1 : _T_131; // @[Mux.scala 47:69]
  assign _T_133 = _T_5[63] ? 6'h0 : _T_132; // @[Mux.scala 47:69]
  assign _GEN_0 = {{63'd0}, _T_5[63:0]}; // @[rawFloatFromIN.scala 55:22]
  assign _T_134 = _GEN_0 << _T_133; // @[rawFloatFromIN.scala 55:22]
  assign _T_140 = {2'h2,~_T_133}; // @[Cat.scala 29:58]
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 72:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 73:23]
  assign roundAnyRawFNToRecFN_io_in_isZero = ~_T_134[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_signedIn & io_in[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(_T_140)}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sig = {{1'd0}, _T_134[63:0]}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[INToRecFN.scala 70:44]
  assign INToRecFN_1_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = INToRecFN_1_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module RecFNToRecFN(
  input  [64:0] io_in,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  RoundAnyRawFNToRecFN_io_invalidExc; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isNaN; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isInf; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isZero; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_sign; // @[RecFNToRecFN.scala 72:19]
  wire [12:0] RoundAnyRawFNToRecFN_io_in_sExp; // @[RecFNToRecFN.scala 72:19]
  wire [53:0] RoundAnyRawFNToRecFN_io_in_sig; // @[RecFNToRecFN.scala 72:19]
  wire [2:0] RoundAnyRawFNToRecFN_io_roundingMode; // @[RecFNToRecFN.scala 72:19]
  wire [32:0] RoundAnyRawFNToRecFN_io_out; // @[RecFNToRecFN.scala 72:19]
  wire [4:0] RoundAnyRawFNToRecFN_io_exceptionFlags; // @[RecFNToRecFN.scala 72:19]
  wire [29:0] RoundAnyRawFNToRecFN_io_covSum; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_metaAssert; // @[RecFNToRecFN.scala 72:19]
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire [1:0] _T_14; // @[Cat.scala 29:58]
  wire [53:0] rawIn_sig; // @[Cat.scala 29:58]
  wire [29:0] RecFNToRecFN_covSum;
  wire [29:0] RoundAnyRawFNToRecFN_sum;
  wire  RoundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_3 RoundAnyRawFNToRecFN ( // @[RecFNToRecFN.scala 72:19]
    .io_invalidExc(RoundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(RoundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(RoundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(RoundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(RoundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(RoundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(RoundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(RoundAnyRawFNToRecFN_io_roundingMode),
    .io_out(RoundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(RoundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(RoundAnyRawFNToRecFN_io_covSum),
    .metaAssert(RoundAnyRawFNToRecFN_metaAssert)
  );
  assign rawIn_isZero = io_in[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_in[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawIn_isNaN = _T_4 & io_in[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign _T_14 = {1'h0,~rawIn_isZero}; // @[Cat.scala 29:58]
  assign rawIn_sig = {1'h0,~rawIn_isZero,io_in[51:0]}; // @[Cat.scala 29:58]
  assign io_out = RoundAnyRawFNToRecFN_io_out; // @[RecFNToRecFN.scala 85:27]
  assign io_exceptionFlags = RoundAnyRawFNToRecFN_io_exceptionFlags; // @[RecFNToRecFN.scala 86:27]
  assign RoundAnyRawFNToRecFN_io_invalidExc = rawIn_isNaN & ~rawIn_sig[51]; // @[RecFNToRecFN.scala 80:48]
  assign RoundAnyRawFNToRecFN_io_in_isNaN = _T_4 & io_in[61]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_isInf = _T_4 & ~io_in[61]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_isZero = io_in[63:61] == 3'h0; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sign = io_in[64]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(io_in[63:52])}; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sig = {_T_14,io_in[51:0]}; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RecFNToRecFN.scala 83:48]
  assign RecFNToRecFN_covSum = 30'h0;
  assign RoundAnyRawFNToRecFN_sum = RecFNToRecFN_covSum + RoundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = RoundAnyRawFNToRecFN_sum;
  assign RoundAnyRawFNToRecFN_metaAssert_wire = RoundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = RoundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module MulAddRecFNPipe_1(
  input         clock,
  input         reset,
  input         io_validin,
  input  [1:0]  io_op,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [64:0] io_c,
  input  [2:0]  io_roundingMode,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output        io_validout,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [1:0] mulAddRecFNToRaw_preMul_io_op; // @[FPU.scala 600:41]
  wire [64:0] mulAddRecFNToRaw_preMul_io_a; // @[FPU.scala 600:41]
  wire [64:0] mulAddRecFNToRaw_preMul_io_b; // @[FPU.scala 600:41]
  wire [64:0] mulAddRecFNToRaw_preMul_io_c; // @[FPU.scala 600:41]
  wire [52:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[FPU.scala 600:41]
  wire [52:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[FPU.scala 600:41]
  wire [105:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FPU.scala 600:41]
  wire [12:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FPU.scala 600:41]
  wire [5:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FPU.scala 600:41]
  wire [54:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FPU.scala 600:41]
  wire [29:0] mulAddRecFNToRaw_preMul_io_covSum; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_preMul_metaAssert; // @[FPU.scala 600:41]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[FPU.scala 601:42]
  wire [12:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[FPU.scala 601:42]
  wire [5:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[FPU.scala 601:42]
  wire [54:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[FPU.scala 601:42]
  wire [106:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[FPU.scala 601:42]
  wire [2:0] mulAddRecFNToRaw_postMul_io_roundingMode; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FPU.scala 601:42]
  wire [12:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FPU.scala 601:42]
  wire [55:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FPU.scala 601:42]
  wire [29:0] mulAddRecFNToRaw_postMul_io_covSum; // @[FPU.scala 601:42]
  wire  mulAddRecFNToRaw_postMul_metaAssert; // @[FPU.scala 601:42]
  wire  roundRawFNToRecFN_io_invalidExc; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_io_in_isInf; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_io_in_isZero; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_io_in_sign; // @[FPU.scala 628:35]
  wire [12:0] roundRawFNToRecFN_io_in_sExp; // @[FPU.scala 628:35]
  wire [55:0] roundRawFNToRecFN_io_in_sig; // @[FPU.scala 628:35]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_io_detectTininess; // @[FPU.scala 628:35]
  wire [64:0] roundRawFNToRecFN_io_out; // @[FPU.scala 628:35]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[FPU.scala 628:35]
  wire [29:0] roundRawFNToRecFN_io_covSum; // @[FPU.scala 628:35]
  wire  roundRawFNToRecFN_metaAssert; // @[FPU.scala 628:35]
  wire [105:0] _T; // @[FPU.scala 609:45]
  wire [106:0] mulAddResult; // @[FPU.scala 610:50]
  reg  _T_2_isSigNaNAny; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg  _T_2_isNaNAOrB; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  _T_2_isInfA; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg  _T_2_isZeroA; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg  _T_2_isInfB; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  _T_2_isZeroB; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  _T_2_signProd; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  _T_2_isNaNC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg  _T_2_isInfC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg  _T_2_isZeroC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [12:0] _T_2_sExpSum; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg  _T_2_doSubMags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg  _T_2_CIsDominant; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [5:0] _T_2_CDom_CAlignDist; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [54:0] _T_2_highAlignedSigC; // @[Reg.scala 15:16]
  reg [63:0] _RAND_14;
  reg  _T_2_bit0AlignedSigC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [106:0] _T_5; // @[Reg.scala 15:16]
  reg [127:0] _RAND_16;
  reg [2:0] _T_8; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [2:0] roundingMode_stage0; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg  detectTininess_stage0; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg  valid_stage0; // @[Valid.scala 117:22]
  reg [31:0] _RAND_20;
  reg  _T_20; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg  _T_23_isNaN; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg  _T_23_isInf; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg  _T_23_isZero; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg  _T_23_sign; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [12:0] _T_23_sExp; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [55:0] _T_23_sig; // @[Reg.scala 15:16]
  reg [63:0] _RAND_27;
  reg [2:0] _T_26; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg  _T_29; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg  _T_31; // @[Valid.scala 117:22]
  reg [31:0] _RAND_30;
  reg  MulAddRecFNPipe_1_state; // @[Register tracking MulAddRecFNPipe_1 state]
  reg [31:0] _RAND_31;
  reg  MulAddRecFNPipe_1_cov [0:1]; // @[Coverage map for MulAddRecFNPipe_1]
  reg [31:0] _RAND_32;
  wire  MulAddRecFNPipe_1_cov_read_data; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_read_addr; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_write_data; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_write_addr; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_write_mask; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_write_en; // @[Coverage map for MulAddRecFNPipe_1]
  reg [29:0] MulAddRecFNPipe_1_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_33;
  wire  valid_stage0_shl;
  wire  valid_stage0_pad;
  wire [29:0] mulAddRecFNToRaw_preMul_sum;
  wire [29:0] mulAddRecFNToRaw_postMul_sum;
  wire [29:0] roundRawFNToRecFN_sum;
  wire  mulAddRecFNToRaw_preMul_metaAssert_wire;
  wire  mulAddRecFNToRaw_postMul_metaAssert_wire;
  wire  roundRawFNToRecFN_metaAssert_wire;
  wire  MulAddRecFNPipe_1_or2;
  wire  MulAddRecFNPipe_1_or0;
  reg  MulAddRecFNPipe_1_metaAssert;
  reg [31:0] _RAND_34;
  MulAddRecFNToRaw_preMul_1 mulAddRecFNToRaw_preMul ( // @[FPU.scala 600:41]
    .io_op(mulAddRecFNToRaw_preMul_io_op),
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC),
    .io_covSum(mulAddRecFNToRaw_preMul_io_covSum),
    .metaAssert(mulAddRecFNToRaw_preMul_metaAssert)
  );
  MulAddRecFNToRaw_postMul_1 mulAddRecFNToRaw_postMul ( // @[FPU.scala 601:42]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_roundingMode(mulAddRecFNToRaw_postMul_io_roundingMode),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig),
    .io_covSum(mulAddRecFNToRaw_postMul_io_covSum),
    .metaAssert(mulAddRecFNToRaw_postMul_metaAssert)
  );
  RoundRawFNToRecFN_3 roundRawFNToRecFN ( // @[FPU.scala 628:35]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundRawFNToRecFN_io_covSum),
    .metaAssert(roundRawFNToRecFN_metaAssert)
  );
  assign _T = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB; // @[FPU.scala 609:45]
  assign mulAddResult = _T + mulAddRecFNToRaw_preMul_io_mulAddC; // @[FPU.scala 610:50]
  assign io_out = roundRawFNToRecFN_io_out; // @[FPU.scala 639:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[FPU.scala 640:23]
  assign io_validout = _T_31; // @[FPU.scala 635:45]
  assign mulAddRecFNToRaw_preMul_io_op = io_op; // @[FPU.scala 603:35]
  assign mulAddRecFNToRaw_preMul_io_a = io_a; // @[FPU.scala 604:35]
  assign mulAddRecFNToRaw_preMul_io_b = io_b; // @[FPU.scala 605:35]
  assign mulAddRecFNToRaw_preMul_io_c = io_c; // @[FPU.scala 606:35]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = _T_2_isSigNaNAny; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = _T_2_isNaNAOrB; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = _T_2_isInfA; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = _T_2_isZeroA; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = _T_2_isInfB; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = _T_2_isZeroB; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = _T_2_signProd; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = _T_2_isNaNC; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = _T_2_isInfC; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = _T_2_isZeroC; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = _T_2_sExpSum; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = _T_2_doSubMags; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = _T_2_CIsDominant; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = _T_2_CDom_CAlignDist; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = _T_2_highAlignedSigC; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = _T_2_bit0AlignedSigC; // @[FPU.scala 618:46]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T_5; // @[FPU.scala 619:46]
  assign mulAddRecFNToRaw_postMul_io_roundingMode = _T_8; // @[FPU.scala 620:46]
  assign roundRawFNToRecFN_io_invalidExc = _T_20; // @[FPU.scala 631:45]
  assign roundRawFNToRecFN_io_infiniteExc = 1'h0; // @[FPU.scala 637:38]
  assign roundRawFNToRecFN_io_in_isNaN = _T_23_isNaN; // @[FPU.scala 632:45]
  assign roundRawFNToRecFN_io_in_isInf = _T_23_isInf; // @[FPU.scala 632:45]
  assign roundRawFNToRecFN_io_in_isZero = _T_23_isZero; // @[FPU.scala 632:45]
  assign roundRawFNToRecFN_io_in_sign = _T_23_sign; // @[FPU.scala 632:45]
  assign roundRawFNToRecFN_io_in_sExp = _T_23_sExp; // @[FPU.scala 632:45]
  assign roundRawFNToRecFN_io_in_sig = _T_23_sig; // @[FPU.scala 632:45]
  assign roundRawFNToRecFN_io_roundingMode = _T_26; // @[FPU.scala 633:45]
  assign roundRawFNToRecFN_io_detectTininess = _T_29; // @[FPU.scala 634:45]
  assign MulAddRecFNPipe_1_cov_read_addr = MulAddRecFNPipe_1_state;
  assign MulAddRecFNPipe_1_cov_read_data = MulAddRecFNPipe_1_cov[MulAddRecFNPipe_1_cov_read_addr]; // @[Coverage map for MulAddRecFNPipe_1]
  assign MulAddRecFNPipe_1_cov_write_data = 1'h1;
  assign MulAddRecFNPipe_1_cov_write_addr = MulAddRecFNPipe_1_state;
  assign MulAddRecFNPipe_1_cov_write_mask = 1'h1;
  assign MulAddRecFNPipe_1_cov_write_en = 1'h1;
  assign valid_stage0_shl = valid_stage0;
  assign valid_stage0_pad = valid_stage0_shl;
  assign mulAddRecFNToRaw_preMul_sum = MulAddRecFNPipe_1_covSum + mulAddRecFNToRaw_preMul_io_covSum;
  assign mulAddRecFNToRaw_postMul_sum = mulAddRecFNToRaw_preMul_sum + mulAddRecFNToRaw_postMul_io_covSum;
  assign roundRawFNToRecFN_sum = mulAddRecFNToRaw_postMul_sum + roundRawFNToRecFN_io_covSum;
  assign io_covSum = roundRawFNToRecFN_sum;
  assign mulAddRecFNToRaw_preMul_metaAssert_wire = mulAddRecFNToRaw_preMul_metaAssert;
  assign mulAddRecFNToRaw_postMul_metaAssert_wire = mulAddRecFNToRaw_postMul_metaAssert;
  assign roundRawFNToRecFN_metaAssert_wire = roundRawFNToRecFN_metaAssert;
  assign MulAddRecFNPipe_1_or2 = mulAddRecFNToRaw_postMul_metaAssert_wire | roundRawFNToRecFN_metaAssert_wire;
  assign MulAddRecFNPipe_1_or0 = mulAddRecFNToRaw_preMul_metaAssert_wire | MulAddRecFNPipe_1_or2;
  assign metaAssert = MulAddRecFNPipe_1_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2_isSigNaNAny = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2_isNaNAOrB = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_isInfA = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2_isZeroA = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2_isInfB = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2_isZeroB = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2_signProd = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2_isNaNC = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2_isInfC = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_2_isZeroC = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2_sExpSum = _RAND_10[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2_doSubMags = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2_CIsDominant = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2_CDom_CAlignDist = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {2{`RANDOM}};
  _T_2_highAlignedSigC = _RAND_14[54:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2_bit0AlignedSigC = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {4{`RANDOM}};
  _T_5 = _RAND_16[106:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_8 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  roundingMode_stage0 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  detectTininess_stage0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  valid_stage0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_20 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_23_isNaN = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_23_isInf = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_23_isZero = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_23_sign = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_23_sExp = _RAND_26[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  _T_23_sig = _RAND_27[55:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_26 = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_31 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  MulAddRecFNPipe_1_state = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    MulAddRecFNPipe_1_cov[initvar] = _RAND_32[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  MulAddRecFNPipe_1_covSum = _RAND_33[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  MulAddRecFNPipe_1_metaAssert = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_2_isSigNaNAny <= 1'h0;
    end else if (io_validin) begin
      _T_2_isSigNaNAny <= mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny;
    end
    if (metaReset) begin
      _T_2_isNaNAOrB <= 1'h0;
    end else if (io_validin) begin
      _T_2_isNaNAOrB <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB;
    end
    if (metaReset) begin
      _T_2_isInfA <= 1'h0;
    end else if (io_validin) begin
      _T_2_isInfA <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfA;
    end
    if (metaReset) begin
      _T_2_isZeroA <= 1'h0;
    end else if (io_validin) begin
      _T_2_isZeroA <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA;
    end
    if (metaReset) begin
      _T_2_isInfB <= 1'h0;
    end else if (io_validin) begin
      _T_2_isInfB <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfB;
    end
    if (metaReset) begin
      _T_2_isZeroB <= 1'h0;
    end else if (io_validin) begin
      _T_2_isZeroB <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB;
    end
    if (metaReset) begin
      _T_2_signProd <= 1'h0;
    end else if (io_validin) begin
      _T_2_signProd <= mulAddRecFNToRaw_preMul_io_toPostMul_signProd;
    end
    if (metaReset) begin
      _T_2_isNaNC <= 1'h0;
    end else if (io_validin) begin
      _T_2_isNaNC <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC;
    end
    if (metaReset) begin
      _T_2_isInfC <= 1'h0;
    end else if (io_validin) begin
      _T_2_isInfC <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfC;
    end
    if (metaReset) begin
      _T_2_isZeroC <= 1'h0;
    end else if (io_validin) begin
      _T_2_isZeroC <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC;
    end
    if (metaReset) begin
      _T_2_sExpSum <= 13'h0;
    end else if (io_validin) begin
      _T_2_sExpSum <= mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum;
    end
    if (metaReset) begin
      _T_2_doSubMags <= 1'h0;
    end else if (io_validin) begin
      _T_2_doSubMags <= mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags;
    end
    if (metaReset) begin
      _T_2_CIsDominant <= 1'h0;
    end else if (io_validin) begin
      _T_2_CIsDominant <= mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant;
    end
    if (metaReset) begin
      _T_2_CDom_CAlignDist <= 6'h0;
    end else if (io_validin) begin
      _T_2_CDom_CAlignDist <= mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist;
    end
    if (metaReset) begin
      _T_2_highAlignedSigC <= 55'h0;
    end else if (io_validin) begin
      _T_2_highAlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC;
    end
    if (metaReset) begin
      _T_2_bit0AlignedSigC <= 1'h0;
    end else if (io_validin) begin
      _T_2_bit0AlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC;
    end
    if (metaReset) begin
      _T_5 <= 107'h0;
    end else if (io_validin) begin
      _T_5 <= mulAddResult;
    end
    if (metaReset) begin
      _T_8 <= 3'h0;
    end else if (io_validin) begin
      _T_8 <= io_roundingMode;
    end
    if (metaReset) begin
      roundingMode_stage0 <= 3'h0;
    end else if (io_validin) begin
      roundingMode_stage0 <= io_roundingMode;
    end
    if (metaReset) begin
      detectTininess_stage0 <= 1'h0;
    end else begin
      detectTininess_stage0 <= io_validin | detectTininess_stage0;
    end
    if (metaReset) begin
      valid_stage0 <= 1'h0;
    end else if (reset) begin
      valid_stage0 <= 1'h0;
    end else begin
      valid_stage0 <= io_validin;
    end
    if (metaReset) begin
      _T_20 <= 1'h0;
    end else if (valid_stage0) begin
      _T_20 <= mulAddRecFNToRaw_postMul_io_invalidExc;
    end
    if (metaReset) begin
      _T_23_isNaN <= 1'h0;
    end else if (valid_stage0) begin
      _T_23_isNaN <= mulAddRecFNToRaw_postMul_io_rawOut_isNaN;
    end
    if (metaReset) begin
      _T_23_isInf <= 1'h0;
    end else if (valid_stage0) begin
      _T_23_isInf <= mulAddRecFNToRaw_postMul_io_rawOut_isInf;
    end
    if (metaReset) begin
      _T_23_isZero <= 1'h0;
    end else if (valid_stage0) begin
      _T_23_isZero <= mulAddRecFNToRaw_postMul_io_rawOut_isZero;
    end
    if (metaReset) begin
      _T_23_sign <= 1'h0;
    end else if (valid_stage0) begin
      _T_23_sign <= mulAddRecFNToRaw_postMul_io_rawOut_sign;
    end
    if (metaReset) begin
      _T_23_sExp <= 13'h0;
    end else if (valid_stage0) begin
      _T_23_sExp <= mulAddRecFNToRaw_postMul_io_rawOut_sExp;
    end
    if (metaReset) begin
      _T_23_sig <= 56'h0;
    end else if (valid_stage0) begin
      _T_23_sig <= mulAddRecFNToRaw_postMul_io_rawOut_sig;
    end
    if (metaReset) begin
      _T_26 <= 3'h0;
    end else if (valid_stage0) begin
      _T_26 <= roundingMode_stage0;
    end
    if (metaReset) begin
      _T_29 <= 1'h0;
    end else if (valid_stage0) begin
      _T_29 <= detectTininess_stage0;
    end
    if (metaReset) begin
      _T_31 <= 1'h0;
    end else if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      _T_31 <= valid_stage0;
    end
    MulAddRecFNPipe_1_state <= valid_stage0_pad;
    if (!(MulAddRecFNPipe_1_cov_read_data)) begin
      MulAddRecFNPipe_1_covSum <= MulAddRecFNPipe_1_covSum + 1'h1;
    end
    if (metaReset) begin
      MulAddRecFNPipe_1_metaAssert <= 1'h0;
    end else begin
      MulAddRecFNPipe_1_metaAssert <= MulAddRecFNPipe_1_metaAssert | MulAddRecFNPipe_1_or0;
    end
  end
  always @(posedge clock) begin
    if(MulAddRecFNPipe_1_cov_write_en & MulAddRecFNPipe_1_cov_write_mask) begin
      MulAddRecFNPipe_1_cov[MulAddRecFNPipe_1_cov_write_addr] <= MulAddRecFNPipe_1_cov_write_data; // @[Coverage map for MulAddRecFNPipe_1]
    end
  end
endmodule
module DivSqrtRecFNToRaw_small(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [2:0]  io_roundingMode,
  output        io_rawOutValid_div,
  output        io_rawOutValid_sqrt,
  output [2:0]  io_roundingModeOut,
  output        io_invalidExc,
  output        io_infiniteExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         divSqrtRawFN_halt
);
  wire  divSqrtRawFN_clock; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_reset; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_inReady; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_inValid; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_sqrtOp; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_a_isNaN; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_a_isInf; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_a_isZero; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_a_sign; // @[DivSqrtRecFN_small.scala 416:15]
  wire [9:0] divSqrtRawFN_io_a_sExp; // @[DivSqrtRecFN_small.scala 416:15]
  wire [24:0] divSqrtRawFN_io_a_sig; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_b_isNaN; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_b_isInf; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_b_isZero; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_b_sign; // @[DivSqrtRecFN_small.scala 416:15]
  wire [9:0] divSqrtRawFN_io_b_sExp; // @[DivSqrtRecFN_small.scala 416:15]
  wire [24:0] divSqrtRawFN_io_b_sig; // @[DivSqrtRecFN_small.scala 416:15]
  wire [2:0] divSqrtRawFN_io_roundingMode; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 416:15]
  wire [2:0] divSqrtRawFN_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_invalidExc; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_infiniteExc; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 416:15]
  wire [9:0] divSqrtRawFN_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 416:15]
  wire [26:0] divSqrtRawFN_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 416:15]
  wire [29:0] divSqrtRawFN_io_covSum; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_metaAssert; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_metaReset; // @[DivSqrtRecFN_small.scala 416:15]
  wire  _T_2; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire  _T_19; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_21; // @[rawFloatFromRecFN.scala 52:54]
  wire [1:0] _T_32; // @[Cat.scala 29:58]
  wire [29:0] DivSqrtRecFNToRaw_small_covSum;
  wire [29:0] divSqrtRawFN_sum;
  wire  divSqrtRawFN_metaAssert_wire;
  reg  DivSqrtRecFNToRaw_small_metaAssert;
  reg [31:0] _RAND_0;
  DivSqrtRawFN_small divSqrtRawFN ( // @[DivSqrtRecFN_small.scala 416:15]
    .clock(divSqrtRawFN_clock),
    .reset(divSqrtRawFN_reset),
    .io_inReady(divSqrtRawFN_io_inReady),
    .io_inValid(divSqrtRawFN_io_inValid),
    .io_sqrtOp(divSqrtRawFN_io_sqrtOp),
    .io_a_isNaN(divSqrtRawFN_io_a_isNaN),
    .io_a_isInf(divSqrtRawFN_io_a_isInf),
    .io_a_isZero(divSqrtRawFN_io_a_isZero),
    .io_a_sign(divSqrtRawFN_io_a_sign),
    .io_a_sExp(divSqrtRawFN_io_a_sExp),
    .io_a_sig(divSqrtRawFN_io_a_sig),
    .io_b_isNaN(divSqrtRawFN_io_b_isNaN),
    .io_b_isInf(divSqrtRawFN_io_b_isInf),
    .io_b_isZero(divSqrtRawFN_io_b_isZero),
    .io_b_sign(divSqrtRawFN_io_b_sign),
    .io_b_sExp(divSqrtRawFN_io_b_sExp),
    .io_b_sig(divSqrtRawFN_io_b_sig),
    .io_roundingMode(divSqrtRawFN_io_roundingMode),
    .io_rawOutValid_div(divSqrtRawFN_io_rawOutValid_div),
    .io_rawOutValid_sqrt(divSqrtRawFN_io_rawOutValid_sqrt),
    .io_roundingModeOut(divSqrtRawFN_io_roundingModeOut),
    .io_invalidExc(divSqrtRawFN_io_invalidExc),
    .io_infiniteExc(divSqrtRawFN_io_infiniteExc),
    .io_rawOut_isNaN(divSqrtRawFN_io_rawOut_isNaN),
    .io_rawOut_isInf(divSqrtRawFN_io_rawOut_isInf),
    .io_rawOut_isZero(divSqrtRawFN_io_rawOut_isZero),
    .io_rawOut_sign(divSqrtRawFN_io_rawOut_sign),
    .io_rawOut_sExp(divSqrtRawFN_io_rawOut_sExp),
    .io_rawOut_sig(divSqrtRawFN_io_rawOut_sig),
    .io_covSum(divSqrtRawFN_io_covSum),
    .metaAssert(divSqrtRawFN_metaAssert),
    .metaReset(divSqrtRawFN_metaReset)
  );
  assign _T_2 = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign _T_15 = {1'h0,~_T_2}; // @[Cat.scala 29:58]
  assign _T_19 = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_21 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign _T_32 = {1'h0,~_T_19}; // @[Cat.scala 29:58]
  assign io_inReady = divSqrtRawFN_io_inReady; // @[DivSqrtRecFN_small.scala 418:16]
  assign io_rawOutValid_div = divSqrtRawFN_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 425:25]
  assign io_rawOutValid_sqrt = divSqrtRawFN_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 426:25]
  assign io_roundingModeOut = divSqrtRawFN_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 427:25]
  assign io_invalidExc = divSqrtRawFN_io_invalidExc; // @[DivSqrtRecFN_small.scala 428:25]
  assign io_infiniteExc = divSqrtRawFN_io_infiniteExc; // @[DivSqrtRecFN_small.scala 429:25]
  assign io_rawOut_isNaN = divSqrtRawFN_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_isInf = divSqrtRawFN_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_isZero = divSqrtRawFN_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_sign = divSqrtRawFN_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_sExp = divSqrtRawFN_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_sig = divSqrtRawFN_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 430:25]
  assign divSqrtRawFN_clock = clock;
  assign divSqrtRawFN_reset = reset;
  assign divSqrtRawFN_io_inValid = io_inValid; // @[DivSqrtRecFN_small.scala 419:34]
  assign divSqrtRawFN_io_sqrtOp = io_sqrtOp; // @[DivSqrtRecFN_small.scala 420:34]
  assign divSqrtRawFN_io_a_isNaN = _T_4 & io_a[29]; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN_io_a_isInf = _T_4 & ~io_a[29]; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN_io_a_isZero = io_a[31:29] == 3'h0; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN_io_a_sign = io_a[32]; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN_io_a_sExp = {1'b0,$signed(io_a[31:23])}; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN_io_a_sig = {_T_15,io_a[22:0]}; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN_io_b_isNaN = _T_21 & io_b[29]; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN_io_b_isInf = _T_21 & ~io_b[29]; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN_io_b_isZero = io_b[31:29] == 3'h0; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN_io_b_sign = io_b[32]; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN_io_b_sExp = {1'b0,$signed(io_b[31:23])}; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN_io_b_sig = {_T_32,io_b[22:0]}; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN_io_roundingMode = io_roundingMode; // @[DivSqrtRecFN_small.scala 423:34]
  assign DivSqrtRecFNToRaw_small_covSum = 30'h0;
  assign divSqrtRawFN_sum = DivSqrtRecFNToRaw_small_covSum + divSqrtRawFN_io_covSum;
  assign io_covSum = divSqrtRawFN_sum;
  assign divSqrtRawFN_metaAssert_wire = divSqrtRawFN_metaAssert;
  assign metaAssert = DivSqrtRecFNToRaw_small_metaAssert;
  assign divSqrtRawFN_metaReset = metaReset | divSqrtRawFN_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DivSqrtRecFNToRaw_small_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      DivSqrtRecFNToRaw_small_metaAssert <= 1'h0;
    end else begin
      DivSqrtRecFNToRaw_small_metaAssert <= DivSqrtRecFNToRaw_small_metaAssert | divSqrtRawFN_metaAssert_wire;
    end
  end
endmodule
module RoundRawFNToRecFN_2(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [9:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [26:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [29:0] RoundRawFNToRecFN_2_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_5 roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundAnyRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundAnyRawFNToRecFN_io_detectTininess),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 316:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_infiniteExc = io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 311:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_detectTininess = io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 314:44]
  assign RoundRawFNToRecFN_2_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = RoundRawFNToRecFN_2_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module DivSqrtRecFNToRaw_small_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [2:0]  io_roundingMode,
  output        io_rawOutValid_div,
  output        io_rawOutValid_sqrt,
  output [2:0]  io_roundingModeOut,
  output        io_invalidExc,
  output        io_infiniteExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [12:0] io_rawOut_sExp,
  output [55:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         divSqrtRawFN_halt
);
  wire  divSqrtRawFN_clock; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_reset; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_inReady; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_inValid; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_sqrtOp; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_a_isNaN; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_a_isInf; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_a_isZero; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_a_sign; // @[DivSqrtRecFN_small.scala 416:15]
  wire [12:0] divSqrtRawFN_io_a_sExp; // @[DivSqrtRecFN_small.scala 416:15]
  wire [53:0] divSqrtRawFN_io_a_sig; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_b_isNaN; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_b_isInf; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_b_isZero; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_b_sign; // @[DivSqrtRecFN_small.scala 416:15]
  wire [12:0] divSqrtRawFN_io_b_sExp; // @[DivSqrtRecFN_small.scala 416:15]
  wire [53:0] divSqrtRawFN_io_b_sig; // @[DivSqrtRecFN_small.scala 416:15]
  wire [2:0] divSqrtRawFN_io_roundingMode; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 416:15]
  wire [2:0] divSqrtRawFN_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_invalidExc; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_infiniteExc; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 416:15]
  wire [12:0] divSqrtRawFN_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 416:15]
  wire [55:0] divSqrtRawFN_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 416:15]
  wire [29:0] divSqrtRawFN_io_covSum; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_metaAssert; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN_metaReset; // @[DivSqrtRecFN_small.scala 416:15]
  wire  _T_2; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire  _T_19; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_21; // @[rawFloatFromRecFN.scala 52:54]
  wire [1:0] _T_32; // @[Cat.scala 29:58]
  wire [29:0] DivSqrtRecFNToRaw_small_1_covSum;
  wire [29:0] divSqrtRawFN_sum;
  wire  divSqrtRawFN_metaAssert_wire;
  reg  DivSqrtRecFNToRaw_small_1_metaAssert;
  reg [31:0] _RAND_0;
  DivSqrtRawFN_small_1 divSqrtRawFN ( // @[DivSqrtRecFN_small.scala 416:15]
    .clock(divSqrtRawFN_clock),
    .reset(divSqrtRawFN_reset),
    .io_inReady(divSqrtRawFN_io_inReady),
    .io_inValid(divSqrtRawFN_io_inValid),
    .io_sqrtOp(divSqrtRawFN_io_sqrtOp),
    .io_a_isNaN(divSqrtRawFN_io_a_isNaN),
    .io_a_isInf(divSqrtRawFN_io_a_isInf),
    .io_a_isZero(divSqrtRawFN_io_a_isZero),
    .io_a_sign(divSqrtRawFN_io_a_sign),
    .io_a_sExp(divSqrtRawFN_io_a_sExp),
    .io_a_sig(divSqrtRawFN_io_a_sig),
    .io_b_isNaN(divSqrtRawFN_io_b_isNaN),
    .io_b_isInf(divSqrtRawFN_io_b_isInf),
    .io_b_isZero(divSqrtRawFN_io_b_isZero),
    .io_b_sign(divSqrtRawFN_io_b_sign),
    .io_b_sExp(divSqrtRawFN_io_b_sExp),
    .io_b_sig(divSqrtRawFN_io_b_sig),
    .io_roundingMode(divSqrtRawFN_io_roundingMode),
    .io_rawOutValid_div(divSqrtRawFN_io_rawOutValid_div),
    .io_rawOutValid_sqrt(divSqrtRawFN_io_rawOutValid_sqrt),
    .io_roundingModeOut(divSqrtRawFN_io_roundingModeOut),
    .io_invalidExc(divSqrtRawFN_io_invalidExc),
    .io_infiniteExc(divSqrtRawFN_io_infiniteExc),
    .io_rawOut_isNaN(divSqrtRawFN_io_rawOut_isNaN),
    .io_rawOut_isInf(divSqrtRawFN_io_rawOut_isInf),
    .io_rawOut_isZero(divSqrtRawFN_io_rawOut_isZero),
    .io_rawOut_sign(divSqrtRawFN_io_rawOut_sign),
    .io_rawOut_sExp(divSqrtRawFN_io_rawOut_sExp),
    .io_rawOut_sig(divSqrtRawFN_io_rawOut_sig),
    .io_covSum(divSqrtRawFN_io_covSum),
    .metaAssert(divSqrtRawFN_metaAssert),
    .metaReset(divSqrtRawFN_metaReset)
  );
  assign _T_2 = io_a[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_a[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign _T_15 = {1'h0,~_T_2}; // @[Cat.scala 29:58]
  assign _T_19 = io_b[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_21 = io_b[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign _T_32 = {1'h0,~_T_19}; // @[Cat.scala 29:58]
  assign io_inReady = divSqrtRawFN_io_inReady; // @[DivSqrtRecFN_small.scala 418:16]
  assign io_rawOutValid_div = divSqrtRawFN_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 425:25]
  assign io_rawOutValid_sqrt = divSqrtRawFN_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 426:25]
  assign io_roundingModeOut = divSqrtRawFN_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 427:25]
  assign io_invalidExc = divSqrtRawFN_io_invalidExc; // @[DivSqrtRecFN_small.scala 428:25]
  assign io_infiniteExc = divSqrtRawFN_io_infiniteExc; // @[DivSqrtRecFN_small.scala 429:25]
  assign io_rawOut_isNaN = divSqrtRawFN_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_isInf = divSqrtRawFN_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_isZero = divSqrtRawFN_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_sign = divSqrtRawFN_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_sExp = divSqrtRawFN_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_sig = divSqrtRawFN_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 430:25]
  assign divSqrtRawFN_clock = clock;
  assign divSqrtRawFN_reset = reset;
  assign divSqrtRawFN_io_inValid = io_inValid; // @[DivSqrtRecFN_small.scala 419:34]
  assign divSqrtRawFN_io_sqrtOp = io_sqrtOp; // @[DivSqrtRecFN_small.scala 420:34]
  assign divSqrtRawFN_io_a_isNaN = _T_4 & io_a[61]; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN_io_a_isInf = _T_4 & ~io_a[61]; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN_io_a_isZero = io_a[63:61] == 3'h0; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN_io_a_sign = io_a[64]; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN_io_a_sExp = {1'b0,$signed(io_a[63:52])}; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN_io_a_sig = {_T_15,io_a[51:0]}; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN_io_b_isNaN = _T_21 & io_b[61]; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN_io_b_isInf = _T_21 & ~io_b[61]; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN_io_b_isZero = io_b[63:61] == 3'h0; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN_io_b_sign = io_b[64]; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN_io_b_sExp = {1'b0,$signed(io_b[63:52])}; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN_io_b_sig = {_T_32,io_b[51:0]}; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN_io_roundingMode = io_roundingMode; // @[DivSqrtRecFN_small.scala 423:34]
  assign DivSqrtRecFNToRaw_small_1_covSum = 30'h0;
  assign divSqrtRawFN_sum = DivSqrtRecFNToRaw_small_1_covSum + divSqrtRawFN_io_covSum;
  assign io_covSum = divSqrtRawFN_sum;
  assign divSqrtRawFN_metaAssert_wire = divSqrtRawFN_metaAssert;
  assign metaAssert = DivSqrtRecFNToRaw_small_1_metaAssert;
  assign divSqrtRawFN_metaReset = metaReset | divSqrtRawFN_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DivSqrtRecFNToRaw_small_1_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      DivSqrtRecFNToRaw_small_1_metaAssert <= 1'h0;
    end else begin
      DivSqrtRecFNToRaw_small_1_metaAssert <= DivSqrtRecFNToRaw_small_1_metaAssert | divSqrtRawFN_metaAssert_wire;
    end
  end
endmodule
module RoundRawFNToRecFN_3(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [55:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [12:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [55:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [64:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [29:0] RoundRawFNToRecFN_3_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_6 roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundAnyRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundAnyRawFNToRecFN_io_detectTininess),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 316:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_infiniteExc = io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 311:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_detectTininess = io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 314:44]
  assign RoundRawFNToRecFN_3_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = RoundRawFNToRecFN_3_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module RVCExpander(
  input  [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0]  io_out_rd,
  output [4:0]  io_out_rs1,
  output [4:0]  io_out_rs2,
  output [4:0]  io_out_rs3,
  output        io_rvc,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  _T_3; // @[RVC.scala 54:29]
  wire [6:0] _T_4; // @[RVC.scala 54:20]
  wire [4:0] _T_14; // @[Cat.scala 29:58]
  wire [29:0] _T_18; // @[Cat.scala 29:58]
  wire [7:0] _T_28; // @[Cat.scala 29:58]
  wire [4:0] _T_30; // @[Cat.scala 29:58]
  wire [27:0] _T_36; // @[Cat.scala 29:58]
  wire [6:0] _T_50; // @[Cat.scala 29:58]
  wire [26:0] _T_58; // @[Cat.scala 29:58]
  wire [27:0] _T_78; // @[Cat.scala 29:58]
  wire [26:0] _T_109; // @[Cat.scala 29:58]
  wire [27:0] _T_136; // @[Cat.scala 29:58]
  wire [26:0] _T_167; // @[Cat.scala 29:58]
  wire [27:0] _T_194; // @[Cat.scala 29:58]
  wire [6:0] _T_205; // @[Bitwise.scala 72:12]
  wire [11:0] _T_207; // @[Cat.scala 29:58]
  wire [31:0] _T_213; // @[Cat.scala 29:58]
  wire  _T_221; // @[RVC.scala 78:24]
  wire [6:0] _T_222; // @[RVC.scala 78:20]
  wire [31:0] _T_233; // @[Cat.scala 29:58]
  wire [31:0] _T_249; // @[Cat.scala 29:58]
  wire  _T_260; // @[RVC.scala 91:29]
  wire [6:0] _T_261; // @[RVC.scala 91:20]
  wire [14:0] _T_264; // @[Bitwise.scala 72:12]
  wire [31:0] _T_267; // @[Cat.scala 29:58]
  wire [31:0] _T_271; // @[Cat.scala 29:58]
  wire  _T_279; // @[RVC.scala 93:14]
  wire  _T_281; // @[RVC.scala 93:27]
  wire  _T_282; // @[RVC.scala 93:21]
  wire [6:0] _T_289; // @[RVC.scala 87:20]
  wire [2:0] _T_292; // @[Bitwise.scala 72:12]
  wire [31:0] _T_307; // @[Cat.scala 29:58]
  wire [31:0] _T_314_bits; // @[RVC.scala 93:10]
  wire [4:0] _T_314_rd; // @[RVC.scala 93:10]
  wire [4:0] _T_314_rs2; // @[RVC.scala 93:10]
  wire [4:0] _T_314_rs3; // @[RVC.scala 93:10]
  wire [25:0] _T_325; // @[Cat.scala 29:58]
  wire [30:0] _GEN_0; // @[RVC.scala 100:23]
  wire [30:0] _T_337; // @[RVC.scala 100:23]
  wire [31:0] _T_350; // @[Cat.scala 29:58]
  wire [2:0] _T_353; // @[Cat.scala 29:58]
  wire  _T_354; // @[package.scala 32:86]
  wire [2:0] _T_355; // @[package.scala 32:76]
  wire  _T_356; // @[package.scala 32:86]
  wire [2:0] _T_357; // @[package.scala 32:76]
  wire  _T_358; // @[package.scala 32:86]
  wire [2:0] _T_359; // @[package.scala 32:76]
  wire  _T_360; // @[package.scala 32:86]
  wire [2:0] _T_361; // @[package.scala 32:76]
  wire  _T_362; // @[package.scala 32:86]
  wire [2:0] _T_363; // @[package.scala 32:76]
  wire  _T_364; // @[package.scala 32:86]
  wire [2:0] _T_365; // @[package.scala 32:76]
  wire  _T_366; // @[package.scala 32:86]
  wire [2:0] _T_367; // @[package.scala 32:76]
  wire  _T_369; // @[RVC.scala 104:30]
  wire [30:0] _T_370; // @[RVC.scala 104:22]
  wire [6:0] _T_372; // @[RVC.scala 105:22]
  wire [24:0] _T_382; // @[Cat.scala 29:58]
  wire [30:0] _GEN_1; // @[RVC.scala 106:43]
  wire [30:0] _T_383; // @[RVC.scala 106:43]
  wire  _T_385; // @[package.scala 32:86]
  wire [30:0] _T_386; // @[package.scala 32:76]
  wire  _T_387; // @[package.scala 32:86]
  wire [31:0] _T_388; // @[package.scala 32:76]
  wire  _T_389; // @[package.scala 32:86]
  wire [31:0] _T_390; // @[package.scala 32:76]
  wire [9:0] _T_401; // @[Bitwise.scala 72:12]
  wire [20:0] _T_416; // @[Cat.scala 29:58]
  wire [31:0] _T_479; // @[Cat.scala 29:58]
  wire [4:0] _T_488; // @[Bitwise.scala 72:12]
  wire [12:0] _T_497; // @[Cat.scala 29:58]
  wire [31:0] _T_546; // @[Cat.scala 29:58]
  wire [31:0] _T_613; // @[Cat.scala 29:58]
  wire [6:0] _T_620; // @[RVC.scala 114:23]
  wire [25:0] _T_629; // @[Cat.scala 29:58]
  wire [28:0] _T_645; // @[Cat.scala 29:58]
  wire [27:0] _T_660; // @[Cat.scala 29:58]
  wire [28:0] _T_675; // @[Cat.scala 29:58]
  wire [24:0] _T_685; // @[Cat.scala 29:58]
  wire [24:0] _T_696; // @[Cat.scala 29:58]
  wire [24:0] _T_707; // @[Cat.scala 29:58]
  wire [24:0] _T_709; // @[Cat.scala 29:58]
  wire [24:0] _T_712; // @[RVC.scala 135:33]
  wire  _T_718; // @[RVC.scala 136:27]
  wire [31:0] _T_689_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_716_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_719_bits; // @[RVC.scala 136:22]
  wire [4:0] _T_719_rd; // @[RVC.scala 136:22]
  wire [4:0] _T_719_rs1; // @[RVC.scala 136:22]
  wire [4:0] _T_719_rs2; // @[RVC.scala 136:22]
  wire [4:0] _T_719_rs3; // @[RVC.scala 136:22]
  wire [24:0] _T_725; // @[Cat.scala 29:58]
  wire [24:0] _T_727; // @[Cat.scala 29:58]
  wire [24:0] _T_728; // @[RVC.scala 138:46]
  wire [24:0] _T_731; // @[RVC.scala 139:33]
  wire [31:0] _T_701_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_735_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_738_bits; // @[RVC.scala 140:25]
  wire [4:0] _T_738_rd; // @[RVC.scala 140:25]
  wire [4:0] _T_738_rs1; // @[RVC.scala 140:25]
  wire [31:0] _T_740_bits; // @[RVC.scala 141:10]
  wire [4:0] _T_740_rd; // @[RVC.scala 141:10]
  wire [4:0] _T_740_rs1; // @[RVC.scala 141:10]
  wire [4:0] _T_740_rs2; // @[RVC.scala 141:10]
  wire [4:0] _T_740_rs3; // @[RVC.scala 141:10]
  wire [8:0] _T_744; // @[Cat.scala 29:58]
  wire [28:0] _T_756; // @[Cat.scala 29:58]
  wire [7:0] _T_764; // @[Cat.scala 29:58]
  wire [27:0] _T_776; // @[Cat.scala 29:58]
  wire [28:0] _T_796; // @[Cat.scala 29:58]
  wire [4:0] _T_843; // @[Cat.scala 29:58]
  wire  _T_844; // @[package.scala 32:86]
  wire [31:0] _T_44_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_24_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_845_bits; // @[package.scala 32:76]
  wire [4:0] _T_845_rd; // @[package.scala 32:76]
  wire [4:0] _T_845_rs1; // @[package.scala 32:76]
  wire [4:0] _T_845_rs3; // @[package.scala 32:76]
  wire  _T_846; // @[package.scala 32:86]
  wire [31:0] _T_66_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_847_bits; // @[package.scala 32:76]
  wire [4:0] _T_847_rd; // @[package.scala 32:76]
  wire [4:0] _T_847_rs1; // @[package.scala 32:76]
  wire [4:0] _T_847_rs3; // @[package.scala 32:76]
  wire  _T_848; // @[package.scala 32:86]
  wire [31:0] _T_86_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_849_bits; // @[package.scala 32:76]
  wire [4:0] _T_849_rd; // @[package.scala 32:76]
  wire [4:0] _T_849_rs1; // @[package.scala 32:76]
  wire [4:0] _T_849_rs3; // @[package.scala 32:76]
  wire  _T_850; // @[package.scala 32:86]
  wire [31:0] _T_117_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_851_bits; // @[package.scala 32:76]
  wire [4:0] _T_851_rd; // @[package.scala 32:76]
  wire [4:0] _T_851_rs1; // @[package.scala 32:76]
  wire [4:0] _T_851_rs3; // @[package.scala 32:76]
  wire  _T_852; // @[package.scala 32:86]
  wire [31:0] _T_144_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_853_bits; // @[package.scala 32:76]
  wire [4:0] _T_853_rd; // @[package.scala 32:76]
  wire [4:0] _T_853_rs1; // @[package.scala 32:76]
  wire [4:0] _T_853_rs3; // @[package.scala 32:76]
  wire  _T_854; // @[package.scala 32:86]
  wire [31:0] _T_175_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_855_bits; // @[package.scala 32:76]
  wire [4:0] _T_855_rd; // @[package.scala 32:76]
  wire [4:0] _T_855_rs1; // @[package.scala 32:76]
  wire [4:0] _T_855_rs3; // @[package.scala 32:76]
  wire  _T_856; // @[package.scala 32:86]
  wire [31:0] _T_202_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_857_bits; // @[package.scala 32:76]
  wire [4:0] _T_857_rd; // @[package.scala 32:76]
  wire [4:0] _T_857_rs1; // @[package.scala 32:76]
  wire [4:0] _T_857_rs3; // @[package.scala 32:76]
  wire  _T_858; // @[package.scala 32:86]
  wire [31:0] _T_859_bits; // @[package.scala 32:76]
  wire [4:0] _T_859_rd; // @[package.scala 32:76]
  wire [4:0] _T_859_rs1; // @[package.scala 32:76]
  wire [4:0] _T_859_rs2; // @[package.scala 32:76]
  wire [4:0] _T_859_rs3; // @[package.scala 32:76]
  wire  _T_860; // @[package.scala 32:86]
  wire [31:0] _T_861_bits; // @[package.scala 32:76]
  wire [4:0] _T_861_rd; // @[package.scala 32:76]
  wire [4:0] _T_861_rs1; // @[package.scala 32:76]
  wire [4:0] _T_861_rs2; // @[package.scala 32:76]
  wire [4:0] _T_861_rs3; // @[package.scala 32:76]
  wire  _T_862; // @[package.scala 32:86]
  wire [31:0] _T_863_bits; // @[package.scala 32:76]
  wire [4:0] _T_863_rd; // @[package.scala 32:76]
  wire [4:0] _T_863_rs1; // @[package.scala 32:76]
  wire [4:0] _T_863_rs2; // @[package.scala 32:76]
  wire [4:0] _T_863_rs3; // @[package.scala 32:76]
  wire  _T_864; // @[package.scala 32:86]
  wire [31:0] _T_865_bits; // @[package.scala 32:76]
  wire [4:0] _T_865_rd; // @[package.scala 32:76]
  wire [4:0] _T_865_rs1; // @[package.scala 32:76]
  wire [4:0] _T_865_rs2; // @[package.scala 32:76]
  wire [4:0] _T_865_rs3; // @[package.scala 32:76]
  wire  _T_866; // @[package.scala 32:86]
  wire [31:0] _T_867_bits; // @[package.scala 32:76]
  wire [4:0] _T_867_rd; // @[package.scala 32:76]
  wire [4:0] _T_867_rs1; // @[package.scala 32:76]
  wire [4:0] _T_867_rs2; // @[package.scala 32:76]
  wire [4:0] _T_867_rs3; // @[package.scala 32:76]
  wire  _T_868; // @[package.scala 32:86]
  wire [31:0] _T_869_bits; // @[package.scala 32:76]
  wire [4:0] _T_869_rd; // @[package.scala 32:76]
  wire [4:0] _T_869_rs1; // @[package.scala 32:76]
  wire [4:0] _T_869_rs2; // @[package.scala 32:76]
  wire [4:0] _T_869_rs3; // @[package.scala 32:76]
  wire  _T_870; // @[package.scala 32:86]
  wire [31:0] _T_871_bits; // @[package.scala 32:76]
  wire [4:0] _T_871_rd; // @[package.scala 32:76]
  wire [4:0] _T_871_rs1; // @[package.scala 32:76]
  wire [4:0] _T_871_rs2; // @[package.scala 32:76]
  wire [4:0] _T_871_rs3; // @[package.scala 32:76]
  wire  _T_872; // @[package.scala 32:86]
  wire [31:0] _T_873_bits; // @[package.scala 32:76]
  wire [4:0] _T_873_rd; // @[package.scala 32:76]
  wire [4:0] _T_873_rs1; // @[package.scala 32:76]
  wire [4:0] _T_873_rs2; // @[package.scala 32:76]
  wire [4:0] _T_873_rs3; // @[package.scala 32:76]
  wire  _T_874; // @[package.scala 32:86]
  wire [31:0] _T_634_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_875_bits; // @[package.scala 32:76]
  wire [4:0] _T_875_rd; // @[package.scala 32:76]
  wire [4:0] _T_875_rs1; // @[package.scala 32:76]
  wire [4:0] _T_875_rs2; // @[package.scala 32:76]
  wire [4:0] _T_875_rs3; // @[package.scala 32:76]
  wire  _T_876; // @[package.scala 32:86]
  wire [31:0] _T_649_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_877_bits; // @[package.scala 32:76]
  wire [4:0] _T_877_rd; // @[package.scala 32:76]
  wire [4:0] _T_877_rs1; // @[package.scala 32:76]
  wire [4:0] _T_877_rs2; // @[package.scala 32:76]
  wire [4:0] _T_877_rs3; // @[package.scala 32:76]
  wire  _T_878; // @[package.scala 32:86]
  wire [31:0] _T_664_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_879_bits; // @[package.scala 32:76]
  wire [4:0] _T_879_rd; // @[package.scala 32:76]
  wire [4:0] _T_879_rs1; // @[package.scala 32:76]
  wire [4:0] _T_879_rs2; // @[package.scala 32:76]
  wire [4:0] _T_879_rs3; // @[package.scala 32:76]
  wire  _T_880; // @[package.scala 32:86]
  wire [31:0] _T_679_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_881_bits; // @[package.scala 32:76]
  wire [4:0] _T_881_rd; // @[package.scala 32:76]
  wire [4:0] _T_881_rs1; // @[package.scala 32:76]
  wire [4:0] _T_881_rs2; // @[package.scala 32:76]
  wire [4:0] _T_881_rs3; // @[package.scala 32:76]
  wire  _T_882; // @[package.scala 32:86]
  wire [31:0] _T_883_bits; // @[package.scala 32:76]
  wire [4:0] _T_883_rd; // @[package.scala 32:76]
  wire [4:0] _T_883_rs1; // @[package.scala 32:76]
  wire [4:0] _T_883_rs2; // @[package.scala 32:76]
  wire [4:0] _T_883_rs3; // @[package.scala 32:76]
  wire  _T_884; // @[package.scala 32:86]
  wire [31:0] _T_760_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_885_bits; // @[package.scala 32:76]
  wire [4:0] _T_885_rd; // @[package.scala 32:76]
  wire [4:0] _T_885_rs1; // @[package.scala 32:76]
  wire [4:0] _T_885_rs2; // @[package.scala 32:76]
  wire [4:0] _T_885_rs3; // @[package.scala 32:76]
  wire  _T_886; // @[package.scala 32:86]
  wire [31:0] _T_780_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_887_bits; // @[package.scala 32:76]
  wire [4:0] _T_887_rd; // @[package.scala 32:76]
  wire [4:0] _T_887_rs1; // @[package.scala 32:76]
  wire [4:0] _T_887_rs2; // @[package.scala 32:76]
  wire [4:0] _T_887_rs3; // @[package.scala 32:76]
  wire  _T_888; // @[package.scala 32:86]
  wire [31:0] _T_800_bits; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _T_889_bits; // @[package.scala 32:76]
  wire [4:0] _T_889_rd; // @[package.scala 32:76]
  wire [4:0] _T_889_rs1; // @[package.scala 32:76]
  wire [4:0] _T_889_rs2; // @[package.scala 32:76]
  wire [4:0] _T_889_rs3; // @[package.scala 32:76]
  wire  _T_890; // @[package.scala 32:86]
  wire [31:0] _T_891_bits; // @[package.scala 32:76]
  wire [4:0] _T_891_rd; // @[package.scala 32:76]
  wire [4:0] _T_891_rs1; // @[package.scala 32:76]
  wire [4:0] _T_891_rs2; // @[package.scala 32:76]
  wire [4:0] _T_891_rs3; // @[package.scala 32:76]
  wire  _T_892; // @[package.scala 32:86]
  wire [31:0] _T_893_bits; // @[package.scala 32:76]
  wire [4:0] _T_893_rd; // @[package.scala 32:76]
  wire [4:0] _T_893_rs1; // @[package.scala 32:76]
  wire [4:0] _T_893_rs2; // @[package.scala 32:76]
  wire [4:0] _T_893_rs3; // @[package.scala 32:76]
  wire  _T_894; // @[package.scala 32:86]
  wire [31:0] _T_895_bits; // @[package.scala 32:76]
  wire [4:0] _T_895_rd; // @[package.scala 32:76]
  wire [4:0] _T_895_rs1; // @[package.scala 32:76]
  wire [4:0] _T_895_rs2; // @[package.scala 32:76]
  wire [4:0] _T_895_rs3; // @[package.scala 32:76]
  wire  _T_896; // @[package.scala 32:86]
  wire [31:0] _T_897_bits; // @[package.scala 32:76]
  wire [4:0] _T_897_rd; // @[package.scala 32:76]
  wire [4:0] _T_897_rs1; // @[package.scala 32:76]
  wire [4:0] _T_897_rs2; // @[package.scala 32:76]
  wire [4:0] _T_897_rs3; // @[package.scala 32:76]
  wire  _T_898; // @[package.scala 32:86]
  wire [31:0] _T_899_bits; // @[package.scala 32:76]
  wire [4:0] _T_899_rd; // @[package.scala 32:76]
  wire [4:0] _T_899_rs1; // @[package.scala 32:76]
  wire [4:0] _T_899_rs2; // @[package.scala 32:76]
  wire [4:0] _T_899_rs3; // @[package.scala 32:76]
  wire  _T_900; // @[package.scala 32:86]
  wire [31:0] _T_901_bits; // @[package.scala 32:76]
  wire [4:0] _T_901_rd; // @[package.scala 32:76]
  wire [4:0] _T_901_rs1; // @[package.scala 32:76]
  wire [4:0] _T_901_rs2; // @[package.scala 32:76]
  wire [4:0] _T_901_rs3; // @[package.scala 32:76]
  wire  _T_902; // @[package.scala 32:86]
  wire [31:0] _T_903_bits; // @[package.scala 32:76]
  wire [4:0] _T_903_rd; // @[package.scala 32:76]
  wire [4:0] _T_903_rs1; // @[package.scala 32:76]
  wire [4:0] _T_903_rs2; // @[package.scala 32:76]
  wire [4:0] _T_903_rs3; // @[package.scala 32:76]
  wire  _T_904; // @[package.scala 32:86]
  wire [29:0] RVCExpander_covSum;
  assign _T_3 = |io_in[12:5]; // @[RVC.scala 54:29]
  assign _T_4 = _T_3 ? 7'h13 : 7'h1f; // @[RVC.scala 54:20]
  assign _T_14 = {2'h1,io_in[4:2]}; // @[Cat.scala 29:58]
  assign _T_18 = {io_in[10:7],io_in[12:11],io_in[5],io_in[6],2'h0,5'h2,3'h0,2'h1,io_in[4:2],_T_4}; // @[Cat.scala 29:58]
  assign _T_28 = {io_in[6:5],io_in[12:10],3'h0}; // @[Cat.scala 29:58]
  assign _T_30 = {2'h1,io_in[9:7]}; // @[Cat.scala 29:58]
  assign _T_36 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h7}; // @[Cat.scala 29:58]
  assign _T_50 = {io_in[5],io_in[12:10],io_in[6],2'h0}; // @[Cat.scala 29:58]
  assign _T_58 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 29:58]
  assign _T_78 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 29:58]
  assign _T_109 = {_T_50[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_50[4:0],7'h3f}; // @[Cat.scala 29:58]
  assign _T_136 = {_T_28[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_T_28[4:0],7'h27}; // @[Cat.scala 29:58]
  assign _T_167 = {_T_50[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_50[4:0],7'h23}; // @[Cat.scala 29:58]
  assign _T_194 = {_T_28[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_T_28[4:0],7'h23}; // @[Cat.scala 29:58]
  assign _T_205 = io_in[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  assign _T_207 = {_T_205,io_in[6:2]}; // @[Cat.scala 29:58]
  assign _T_213 = {_T_205,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13}; // @[Cat.scala 29:58]
  assign _T_221 = |io_in[11:7]; // @[RVC.scala 78:24]
  assign _T_222 = _T_221 ? 7'h1b : 7'h1f; // @[RVC.scala 78:20]
  assign _T_233 = {_T_205,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],_T_222}; // @[Cat.scala 29:58]
  assign _T_249 = {_T_205,io_in[6:2],5'h0,3'h0,io_in[11:7],7'h13}; // @[Cat.scala 29:58]
  assign _T_260 = |_T_207; // @[RVC.scala 91:29]
  assign _T_261 = _T_260 ? 7'h37 : 7'h3f; // @[RVC.scala 91:20]
  assign _T_264 = io_in[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  assign _T_267 = {_T_264,io_in[6:2],12'h0}; // @[Cat.scala 29:58]
  assign _T_271 = {_T_267[31:12],io_in[11:7],_T_261}; // @[Cat.scala 29:58]
  assign _T_279 = io_in[11:7] == 5'h0; // @[RVC.scala 93:14]
  assign _T_281 = io_in[11:7] == 5'h2; // @[RVC.scala 93:27]
  assign _T_282 = _T_279 | _T_281; // @[RVC.scala 93:21]
  assign _T_289 = _T_260 ? 7'h13 : 7'h1f; // @[RVC.scala 87:20]
  assign _T_292 = io_in[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  assign _T_307 = {_T_292,io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[11:7],_T_289}; // @[Cat.scala 29:58]
  assign _T_314_bits = _T_282 ? _T_307 : _T_271; // @[RVC.scala 93:10]
  assign _T_314_rd = _T_282 ? io_in[11:7] : io_in[11:7]; // @[RVC.scala 93:10]
  assign _T_314_rs2 = _T_282 ? _T_14 : _T_14; // @[RVC.scala 93:10]
  assign _T_314_rs3 = _T_282 ? io_in[31:27] : io_in[31:27]; // @[RVC.scala 93:10]
  assign _T_325 = {io_in[12],io_in[6:2],2'h1,io_in[9:7],3'h5,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 29:58]
  assign _GEN_0 = {{5'd0}, _T_325}; // @[RVC.scala 100:23]
  assign _T_337 = _GEN_0 | 31'h40000000; // @[RVC.scala 100:23]
  assign _T_350 = {_T_205,io_in[6:2],2'h1,io_in[9:7],3'h7,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 29:58]
  assign _T_353 = {io_in[12],io_in[6:5]}; // @[Cat.scala 29:58]
  assign _T_354 = _T_353 == 3'h1; // @[package.scala 32:86]
  assign _T_355 = _T_354 ? 3'h4 : 3'h0; // @[package.scala 32:76]
  assign _T_356 = _T_353 == 3'h2; // @[package.scala 32:86]
  assign _T_357 = _T_356 ? 3'h6 : _T_355; // @[package.scala 32:76]
  assign _T_358 = _T_353 == 3'h3; // @[package.scala 32:86]
  assign _T_359 = _T_358 ? 3'h7 : _T_357; // @[package.scala 32:76]
  assign _T_360 = _T_353 == 3'h4; // @[package.scala 32:86]
  assign _T_361 = _T_360 ? 3'h0 : _T_359; // @[package.scala 32:76]
  assign _T_362 = _T_353 == 3'h5; // @[package.scala 32:86]
  assign _T_363 = _T_362 ? 3'h0 : _T_361; // @[package.scala 32:76]
  assign _T_364 = _T_353 == 3'h6; // @[package.scala 32:86]
  assign _T_365 = _T_364 ? 3'h2 : _T_363; // @[package.scala 32:76]
  assign _T_366 = _T_353 == 3'h7; // @[package.scala 32:86]
  assign _T_367 = _T_366 ? 3'h3 : _T_365; // @[package.scala 32:76]
  assign _T_369 = io_in[6:5] == 2'h0; // @[RVC.scala 104:30]
  assign _T_370 = _T_369 ? 31'h40000000 : 31'h0; // @[RVC.scala 104:22]
  assign _T_372 = io_in[12] ? 7'h3b : 7'h33; // @[RVC.scala 105:22]
  assign _T_382 = {2'h1,io_in[4:2],2'h1,io_in[9:7],_T_367,2'h1,io_in[9:7],_T_372}; // @[Cat.scala 29:58]
  assign _GEN_1 = {{6'd0}, _T_382}; // @[RVC.scala 106:43]
  assign _T_383 = _GEN_1 | _T_370; // @[RVC.scala 106:43]
  assign _T_385 = io_in[11:10] == 2'h1; // @[package.scala 32:86]
  assign _T_386 = _T_385 ? _T_337 : {{5'd0}, _T_325}; // @[package.scala 32:76]
  assign _T_387 = io_in[11:10] == 2'h2; // @[package.scala 32:86]
  assign _T_388 = _T_387 ? _T_350 : {{1'd0}, _T_386}; // @[package.scala 32:76]
  assign _T_389 = io_in[11:10] == 2'h3; // @[package.scala 32:86]
  assign _T_390 = _T_389 ? {{1'd0}, _T_383} : _T_388; // @[package.scala 32:76]
  assign _T_401 = io_in[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  assign _T_416 = {_T_401,io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],1'h0}; // @[Cat.scala 29:58]
  assign _T_479 = {_T_416[20],_T_416[10:1],_T_416[11],_T_416[19:12],5'h0,7'h6f}; // @[Cat.scala 29:58]
  assign _T_488 = io_in[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  assign _T_497 = {_T_488,io_in[6:5],io_in[2],io_in[11:10],io_in[4:3],1'h0}; // @[Cat.scala 29:58]
  assign _T_546 = {_T_497[12],_T_497[10:5],5'h0,2'h1,io_in[9:7],3'h0,_T_497[4:1],_T_497[11],7'h63}; // @[Cat.scala 29:58]
  assign _T_613 = {_T_497[12],_T_497[10:5],5'h0,2'h1,io_in[9:7],3'h1,_T_497[4:1],_T_497[11],7'h63}; // @[Cat.scala 29:58]
  assign _T_620 = _T_221 ? 7'h3 : 7'h1f; // @[RVC.scala 114:23]
  assign _T_629 = {io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13}; // @[Cat.scala 29:58]
  assign _T_645 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],7'h7}; // @[Cat.scala 29:58]
  assign _T_660 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],_T_620}; // @[Cat.scala 29:58]
  assign _T_675 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],_T_620}; // @[Cat.scala 29:58]
  assign _T_685 = {io_in[6:2],5'h0,3'h0,io_in[11:7],7'h33}; // @[Cat.scala 29:58]
  assign _T_696 = {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33}; // @[Cat.scala 29:58]
  assign _T_707 = {io_in[6:2],io_in[11:7],3'h0,12'h67}; // @[Cat.scala 29:58]
  assign _T_709 = {_T_707[24:7],7'h1f}; // @[Cat.scala 29:58]
  assign _T_712 = _T_221 ? _T_707 : _T_709; // @[RVC.scala 135:33]
  assign _T_718 = |io_in[6:2]; // @[RVC.scala 136:27]
  assign _T_689_bits = {{7'd0}, _T_685}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_716_bits = {{7'd0}, _T_712}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_719_bits = _T_718 ? _T_689_bits : _T_716_bits; // @[RVC.scala 136:22]
  assign _T_719_rd = _T_718 ? io_in[11:7] : 5'h0; // @[RVC.scala 136:22]
  assign _T_719_rs1 = _T_718 ? 5'h0 : io_in[11:7]; // @[RVC.scala 136:22]
  assign _T_719_rs2 = _T_718 ? io_in[6:2] : io_in[6:2]; // @[RVC.scala 136:22]
  assign _T_719_rs3 = _T_718 ? io_in[31:27] : io_in[31:27]; // @[RVC.scala 136:22]
  assign _T_725 = {io_in[6:2],io_in[11:7],3'h0,12'he7}; // @[Cat.scala 29:58]
  assign _T_727 = {_T_707[24:7],7'h73}; // @[Cat.scala 29:58]
  assign _T_728 = _T_727 | 25'h100000; // @[RVC.scala 138:46]
  assign _T_731 = _T_221 ? _T_725 : _T_728; // @[RVC.scala 139:33]
  assign _T_701_bits = {{7'd0}, _T_696}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_735_bits = {{7'd0}, _T_731}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_738_bits = _T_718 ? _T_701_bits : _T_735_bits; // @[RVC.scala 140:25]
  assign _T_738_rd = _T_718 ? io_in[11:7] : 5'h1; // @[RVC.scala 140:25]
  assign _T_738_rs1 = _T_718 ? io_in[11:7] : io_in[11:7]; // @[RVC.scala 140:25]
  assign _T_740_bits = io_in[12] ? _T_738_bits : _T_719_bits; // @[RVC.scala 141:10]
  assign _T_740_rd = io_in[12] ? _T_738_rd : _T_719_rd; // @[RVC.scala 141:10]
  assign _T_740_rs1 = io_in[12] ? _T_738_rs1 : _T_719_rs1; // @[RVC.scala 141:10]
  assign _T_740_rs2 = io_in[12] ? _T_719_rs2 : _T_719_rs2; // @[RVC.scala 141:10]
  assign _T_740_rs3 = io_in[12] ? _T_719_rs3 : _T_719_rs3; // @[RVC.scala 141:10]
  assign _T_744 = {io_in[9:7],io_in[12:10],3'h0}; // @[Cat.scala 29:58]
  assign _T_756 = {_T_744[8:5],io_in[6:2],5'h2,3'h3,_T_744[4:0],7'h27}; // @[Cat.scala 29:58]
  assign _T_764 = {io_in[8:7],io_in[12:9],2'h0}; // @[Cat.scala 29:58]
  assign _T_776 = {_T_764[7:5],io_in[6:2],5'h2,3'h2,_T_764[4:0],7'h23}; // @[Cat.scala 29:58]
  assign _T_796 = {_T_744[8:5],io_in[6:2],5'h2,3'h3,_T_744[4:0],7'h23}; // @[Cat.scala 29:58]
  assign _T_843 = {io_in[1:0],io_in[15:13]}; // @[Cat.scala 29:58]
  assign _T_844 = _T_843 == 5'h1; // @[package.scala 32:86]
  assign _T_44_bits = {{4'd0}, _T_36}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_24_bits = {{2'd0}, _T_18}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_845_bits = _T_844 ? _T_44_bits : _T_24_bits; // @[package.scala 32:76]
  assign _T_845_rd = _T_844 ? _T_14 : _T_14; // @[package.scala 32:76]
  assign _T_845_rs1 = _T_844 ? _T_30 : 5'h2; // @[package.scala 32:76]
  assign _T_845_rs3 = _T_844 ? io_in[31:27] : io_in[31:27]; // @[package.scala 32:76]
  assign _T_846 = _T_843 == 5'h2; // @[package.scala 32:86]
  assign _T_66_bits = {{5'd0}, _T_58}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_847_bits = _T_846 ? _T_66_bits : _T_845_bits; // @[package.scala 32:76]
  assign _T_847_rd = _T_846 ? _T_14 : _T_845_rd; // @[package.scala 32:76]
  assign _T_847_rs1 = _T_846 ? _T_30 : _T_845_rs1; // @[package.scala 32:76]
  assign _T_847_rs3 = _T_846 ? io_in[31:27] : _T_845_rs3; // @[package.scala 32:76]
  assign _T_848 = _T_843 == 5'h3; // @[package.scala 32:86]
  assign _T_86_bits = {{4'd0}, _T_78}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_849_bits = _T_848 ? _T_86_bits : _T_847_bits; // @[package.scala 32:76]
  assign _T_849_rd = _T_848 ? _T_14 : _T_847_rd; // @[package.scala 32:76]
  assign _T_849_rs1 = _T_848 ? _T_30 : _T_847_rs1; // @[package.scala 32:76]
  assign _T_849_rs3 = _T_848 ? io_in[31:27] : _T_847_rs3; // @[package.scala 32:76]
  assign _T_850 = _T_843 == 5'h4; // @[package.scala 32:86]
  assign _T_117_bits = {{5'd0}, _T_109}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_851_bits = _T_850 ? _T_117_bits : _T_849_bits; // @[package.scala 32:76]
  assign _T_851_rd = _T_850 ? _T_14 : _T_849_rd; // @[package.scala 32:76]
  assign _T_851_rs1 = _T_850 ? _T_30 : _T_849_rs1; // @[package.scala 32:76]
  assign _T_851_rs3 = _T_850 ? io_in[31:27] : _T_849_rs3; // @[package.scala 32:76]
  assign _T_852 = _T_843 == 5'h5; // @[package.scala 32:86]
  assign _T_144_bits = {{4'd0}, _T_136}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_853_bits = _T_852 ? _T_144_bits : _T_851_bits; // @[package.scala 32:76]
  assign _T_853_rd = _T_852 ? _T_14 : _T_851_rd; // @[package.scala 32:76]
  assign _T_853_rs1 = _T_852 ? _T_30 : _T_851_rs1; // @[package.scala 32:76]
  assign _T_853_rs3 = _T_852 ? io_in[31:27] : _T_851_rs3; // @[package.scala 32:76]
  assign _T_854 = _T_843 == 5'h6; // @[package.scala 32:86]
  assign _T_175_bits = {{5'd0}, _T_167}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_855_bits = _T_854 ? _T_175_bits : _T_853_bits; // @[package.scala 32:76]
  assign _T_855_rd = _T_854 ? _T_14 : _T_853_rd; // @[package.scala 32:76]
  assign _T_855_rs1 = _T_854 ? _T_30 : _T_853_rs1; // @[package.scala 32:76]
  assign _T_855_rs3 = _T_854 ? io_in[31:27] : _T_853_rs3; // @[package.scala 32:76]
  assign _T_856 = _T_843 == 5'h7; // @[package.scala 32:86]
  assign _T_202_bits = {{4'd0}, _T_194}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_857_bits = _T_856 ? _T_202_bits : _T_855_bits; // @[package.scala 32:76]
  assign _T_857_rd = _T_856 ? _T_14 : _T_855_rd; // @[package.scala 32:76]
  assign _T_857_rs1 = _T_856 ? _T_30 : _T_855_rs1; // @[package.scala 32:76]
  assign _T_857_rs3 = _T_856 ? io_in[31:27] : _T_855_rs3; // @[package.scala 32:76]
  assign _T_858 = _T_843 == 5'h8; // @[package.scala 32:86]
  assign _T_859_bits = _T_858 ? _T_213 : _T_857_bits; // @[package.scala 32:76]
  assign _T_859_rd = _T_858 ? io_in[11:7] : _T_857_rd; // @[package.scala 32:76]
  assign _T_859_rs1 = _T_858 ? io_in[11:7] : _T_857_rs1; // @[package.scala 32:76]
  assign _T_859_rs2 = _T_858 ? _T_14 : _T_857_rd; // @[package.scala 32:76]
  assign _T_859_rs3 = _T_858 ? io_in[31:27] : _T_857_rs3; // @[package.scala 32:76]
  assign _T_860 = _T_843 == 5'h9; // @[package.scala 32:86]
  assign _T_861_bits = _T_860 ? _T_233 : _T_859_bits; // @[package.scala 32:76]
  assign _T_861_rd = _T_860 ? io_in[11:7] : _T_859_rd; // @[package.scala 32:76]
  assign _T_861_rs1 = _T_860 ? io_in[11:7] : _T_859_rs1; // @[package.scala 32:76]
  assign _T_861_rs2 = _T_860 ? _T_14 : _T_859_rs2; // @[package.scala 32:76]
  assign _T_861_rs3 = _T_860 ? io_in[31:27] : _T_859_rs3; // @[package.scala 32:76]
  assign _T_862 = _T_843 == 5'ha; // @[package.scala 32:86]
  assign _T_863_bits = _T_862 ? _T_249 : _T_861_bits; // @[package.scala 32:76]
  assign _T_863_rd = _T_862 ? io_in[11:7] : _T_861_rd; // @[package.scala 32:76]
  assign _T_863_rs1 = _T_862 ? 5'h0 : _T_861_rs1; // @[package.scala 32:76]
  assign _T_863_rs2 = _T_862 ? _T_14 : _T_861_rs2; // @[package.scala 32:76]
  assign _T_863_rs3 = _T_862 ? io_in[31:27] : _T_861_rs3; // @[package.scala 32:76]
  assign _T_864 = _T_843 == 5'hb; // @[package.scala 32:86]
  assign _T_865_bits = _T_864 ? _T_314_bits : _T_863_bits; // @[package.scala 32:76]
  assign _T_865_rd = _T_864 ? _T_314_rd : _T_863_rd; // @[package.scala 32:76]
  assign _T_865_rs1 = _T_864 ? _T_314_rd : _T_863_rs1; // @[package.scala 32:76]
  assign _T_865_rs2 = _T_864 ? _T_314_rs2 : _T_863_rs2; // @[package.scala 32:76]
  assign _T_865_rs3 = _T_864 ? _T_314_rs3 : _T_863_rs3; // @[package.scala 32:76]
  assign _T_866 = _T_843 == 5'hc; // @[package.scala 32:86]
  assign _T_867_bits = _T_866 ? _T_390 : _T_865_bits; // @[package.scala 32:76]
  assign _T_867_rd = _T_866 ? _T_30 : _T_865_rd; // @[package.scala 32:76]
  assign _T_867_rs1 = _T_866 ? _T_30 : _T_865_rs1; // @[package.scala 32:76]
  assign _T_867_rs2 = _T_866 ? _T_14 : _T_865_rs2; // @[package.scala 32:76]
  assign _T_867_rs3 = _T_866 ? io_in[31:27] : _T_865_rs3; // @[package.scala 32:76]
  assign _T_868 = _T_843 == 5'hd; // @[package.scala 32:86]
  assign _T_869_bits = _T_868 ? _T_479 : _T_867_bits; // @[package.scala 32:76]
  assign _T_869_rd = _T_868 ? 5'h0 : _T_867_rd; // @[package.scala 32:76]
  assign _T_869_rs1 = _T_868 ? _T_30 : _T_867_rs1; // @[package.scala 32:76]
  assign _T_869_rs2 = _T_868 ? _T_14 : _T_867_rs2; // @[package.scala 32:76]
  assign _T_869_rs3 = _T_868 ? io_in[31:27] : _T_867_rs3; // @[package.scala 32:76]
  assign _T_870 = _T_843 == 5'he; // @[package.scala 32:86]
  assign _T_871_bits = _T_870 ? _T_546 : _T_869_bits; // @[package.scala 32:76]
  assign _T_871_rd = _T_870 ? _T_30 : _T_869_rd; // @[package.scala 32:76]
  assign _T_871_rs1 = _T_870 ? _T_30 : _T_869_rs1; // @[package.scala 32:76]
  assign _T_871_rs2 = _T_870 ? 5'h0 : _T_869_rs2; // @[package.scala 32:76]
  assign _T_871_rs3 = _T_870 ? io_in[31:27] : _T_869_rs3; // @[package.scala 32:76]
  assign _T_872 = _T_843 == 5'hf; // @[package.scala 32:86]
  assign _T_873_bits = _T_872 ? _T_613 : _T_871_bits; // @[package.scala 32:76]
  assign _T_873_rd = _T_872 ? 5'h0 : _T_871_rd; // @[package.scala 32:76]
  assign _T_873_rs1 = _T_872 ? _T_30 : _T_871_rs1; // @[package.scala 32:76]
  assign _T_873_rs2 = _T_872 ? 5'h0 : _T_871_rs2; // @[package.scala 32:76]
  assign _T_873_rs3 = _T_872 ? io_in[31:27] : _T_871_rs3; // @[package.scala 32:76]
  assign _T_874 = _T_843 == 5'h10; // @[package.scala 32:86]
  assign _T_634_bits = {{6'd0}, _T_629}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_875_bits = _T_874 ? _T_634_bits : _T_873_bits; // @[package.scala 32:76]
  assign _T_875_rd = _T_874 ? io_in[11:7] : _T_873_rd; // @[package.scala 32:76]
  assign _T_875_rs1 = _T_874 ? io_in[11:7] : _T_873_rs1; // @[package.scala 32:76]
  assign _T_875_rs2 = _T_874 ? io_in[6:2] : _T_873_rs2; // @[package.scala 32:76]
  assign _T_875_rs3 = _T_874 ? io_in[31:27] : _T_873_rs3; // @[package.scala 32:76]
  assign _T_876 = _T_843 == 5'h11; // @[package.scala 32:86]
  assign _T_649_bits = {{3'd0}, _T_645}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_877_bits = _T_876 ? _T_649_bits : _T_875_bits; // @[package.scala 32:76]
  assign _T_877_rd = _T_876 ? io_in[11:7] : _T_875_rd; // @[package.scala 32:76]
  assign _T_877_rs1 = _T_876 ? 5'h2 : _T_875_rs1; // @[package.scala 32:76]
  assign _T_877_rs2 = _T_876 ? io_in[6:2] : _T_875_rs2; // @[package.scala 32:76]
  assign _T_877_rs3 = _T_876 ? io_in[31:27] : _T_875_rs3; // @[package.scala 32:76]
  assign _T_878 = _T_843 == 5'h12; // @[package.scala 32:86]
  assign _T_664_bits = {{4'd0}, _T_660}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_879_bits = _T_878 ? _T_664_bits : _T_877_bits; // @[package.scala 32:76]
  assign _T_879_rd = _T_878 ? io_in[11:7] : _T_877_rd; // @[package.scala 32:76]
  assign _T_879_rs1 = _T_878 ? 5'h2 : _T_877_rs1; // @[package.scala 32:76]
  assign _T_879_rs2 = _T_878 ? io_in[6:2] : _T_877_rs2; // @[package.scala 32:76]
  assign _T_879_rs3 = _T_878 ? io_in[31:27] : _T_877_rs3; // @[package.scala 32:76]
  assign _T_880 = _T_843 == 5'h13; // @[package.scala 32:86]
  assign _T_679_bits = {{3'd0}, _T_675}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_881_bits = _T_880 ? _T_679_bits : _T_879_bits; // @[package.scala 32:76]
  assign _T_881_rd = _T_880 ? io_in[11:7] : _T_879_rd; // @[package.scala 32:76]
  assign _T_881_rs1 = _T_880 ? 5'h2 : _T_879_rs1; // @[package.scala 32:76]
  assign _T_881_rs2 = _T_880 ? io_in[6:2] : _T_879_rs2; // @[package.scala 32:76]
  assign _T_881_rs3 = _T_880 ? io_in[31:27] : _T_879_rs3; // @[package.scala 32:76]
  assign _T_882 = _T_843 == 5'h14; // @[package.scala 32:86]
  assign _T_883_bits = _T_882 ? _T_740_bits : _T_881_bits; // @[package.scala 32:76]
  assign _T_883_rd = _T_882 ? _T_740_rd : _T_881_rd; // @[package.scala 32:76]
  assign _T_883_rs1 = _T_882 ? _T_740_rs1 : _T_881_rs1; // @[package.scala 32:76]
  assign _T_883_rs2 = _T_882 ? _T_740_rs2 : _T_881_rs2; // @[package.scala 32:76]
  assign _T_883_rs3 = _T_882 ? _T_740_rs3 : _T_881_rs3; // @[package.scala 32:76]
  assign _T_884 = _T_843 == 5'h15; // @[package.scala 32:86]
  assign _T_760_bits = {{3'd0}, _T_756}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_885_bits = _T_884 ? _T_760_bits : _T_883_bits; // @[package.scala 32:76]
  assign _T_885_rd = _T_884 ? io_in[11:7] : _T_883_rd; // @[package.scala 32:76]
  assign _T_885_rs1 = _T_884 ? 5'h2 : _T_883_rs1; // @[package.scala 32:76]
  assign _T_885_rs2 = _T_884 ? io_in[6:2] : _T_883_rs2; // @[package.scala 32:76]
  assign _T_885_rs3 = _T_884 ? io_in[31:27] : _T_883_rs3; // @[package.scala 32:76]
  assign _T_886 = _T_843 == 5'h16; // @[package.scala 32:86]
  assign _T_780_bits = {{4'd0}, _T_776}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_887_bits = _T_886 ? _T_780_bits : _T_885_bits; // @[package.scala 32:76]
  assign _T_887_rd = _T_886 ? io_in[11:7] : _T_885_rd; // @[package.scala 32:76]
  assign _T_887_rs1 = _T_886 ? 5'h2 : _T_885_rs1; // @[package.scala 32:76]
  assign _T_887_rs2 = _T_886 ? io_in[6:2] : _T_885_rs2; // @[package.scala 32:76]
  assign _T_887_rs3 = _T_886 ? io_in[31:27] : _T_885_rs3; // @[package.scala 32:76]
  assign _T_888 = _T_843 == 5'h17; // @[package.scala 32:86]
  assign _T_800_bits = {{3'd0}, _T_796}; // @[RVC.scala 22:19 RVC.scala 23:14]
  assign _T_889_bits = _T_888 ? _T_800_bits : _T_887_bits; // @[package.scala 32:76]
  assign _T_889_rd = _T_888 ? io_in[11:7] : _T_887_rd; // @[package.scala 32:76]
  assign _T_889_rs1 = _T_888 ? 5'h2 : _T_887_rs1; // @[package.scala 32:76]
  assign _T_889_rs2 = _T_888 ? io_in[6:2] : _T_887_rs2; // @[package.scala 32:76]
  assign _T_889_rs3 = _T_888 ? io_in[31:27] : _T_887_rs3; // @[package.scala 32:76]
  assign _T_890 = _T_843 == 5'h18; // @[package.scala 32:86]
  assign _T_891_bits = _T_890 ? io_in : _T_889_bits; // @[package.scala 32:76]
  assign _T_891_rd = _T_890 ? io_in[11:7] : _T_889_rd; // @[package.scala 32:76]
  assign _T_891_rs1 = _T_890 ? io_in[19:15] : _T_889_rs1; // @[package.scala 32:76]
  assign _T_891_rs2 = _T_890 ? io_in[24:20] : _T_889_rs2; // @[package.scala 32:76]
  assign _T_891_rs3 = _T_890 ? io_in[31:27] : _T_889_rs3; // @[package.scala 32:76]
  assign _T_892 = _T_843 == 5'h19; // @[package.scala 32:86]
  assign _T_893_bits = _T_892 ? io_in : _T_891_bits; // @[package.scala 32:76]
  assign _T_893_rd = _T_892 ? io_in[11:7] : _T_891_rd; // @[package.scala 32:76]
  assign _T_893_rs1 = _T_892 ? io_in[19:15] : _T_891_rs1; // @[package.scala 32:76]
  assign _T_893_rs2 = _T_892 ? io_in[24:20] : _T_891_rs2; // @[package.scala 32:76]
  assign _T_893_rs3 = _T_892 ? io_in[31:27] : _T_891_rs3; // @[package.scala 32:76]
  assign _T_894 = _T_843 == 5'h1a; // @[package.scala 32:86]
  assign _T_895_bits = _T_894 ? io_in : _T_893_bits; // @[package.scala 32:76]
  assign _T_895_rd = _T_894 ? io_in[11:7] : _T_893_rd; // @[package.scala 32:76]
  assign _T_895_rs1 = _T_894 ? io_in[19:15] : _T_893_rs1; // @[package.scala 32:76]
  assign _T_895_rs2 = _T_894 ? io_in[24:20] : _T_893_rs2; // @[package.scala 32:76]
  assign _T_895_rs3 = _T_894 ? io_in[31:27] : _T_893_rs3; // @[package.scala 32:76]
  assign _T_896 = _T_843 == 5'h1b; // @[package.scala 32:86]
  assign _T_897_bits = _T_896 ? io_in : _T_895_bits; // @[package.scala 32:76]
  assign _T_897_rd = _T_896 ? io_in[11:7] : _T_895_rd; // @[package.scala 32:76]
  assign _T_897_rs1 = _T_896 ? io_in[19:15] : _T_895_rs1; // @[package.scala 32:76]
  assign _T_897_rs2 = _T_896 ? io_in[24:20] : _T_895_rs2; // @[package.scala 32:76]
  assign _T_897_rs3 = _T_896 ? io_in[31:27] : _T_895_rs3; // @[package.scala 32:76]
  assign _T_898 = _T_843 == 5'h1c; // @[package.scala 32:86]
  assign _T_899_bits = _T_898 ? io_in : _T_897_bits; // @[package.scala 32:76]
  assign _T_899_rd = _T_898 ? io_in[11:7] : _T_897_rd; // @[package.scala 32:76]
  assign _T_899_rs1 = _T_898 ? io_in[19:15] : _T_897_rs1; // @[package.scala 32:76]
  assign _T_899_rs2 = _T_898 ? io_in[24:20] : _T_897_rs2; // @[package.scala 32:76]
  assign _T_899_rs3 = _T_898 ? io_in[31:27] : _T_897_rs3; // @[package.scala 32:76]
  assign _T_900 = _T_843 == 5'h1d; // @[package.scala 32:86]
  assign _T_901_bits = _T_900 ? io_in : _T_899_bits; // @[package.scala 32:76]
  assign _T_901_rd = _T_900 ? io_in[11:7] : _T_899_rd; // @[package.scala 32:76]
  assign _T_901_rs1 = _T_900 ? io_in[19:15] : _T_899_rs1; // @[package.scala 32:76]
  assign _T_901_rs2 = _T_900 ? io_in[24:20] : _T_899_rs2; // @[package.scala 32:76]
  assign _T_901_rs3 = _T_900 ? io_in[31:27] : _T_899_rs3; // @[package.scala 32:76]
  assign _T_902 = _T_843 == 5'h1e; // @[package.scala 32:86]
  assign _T_903_bits = _T_902 ? io_in : _T_901_bits; // @[package.scala 32:76]
  assign _T_903_rd = _T_902 ? io_in[11:7] : _T_901_rd; // @[package.scala 32:76]
  assign _T_903_rs1 = _T_902 ? io_in[19:15] : _T_901_rs1; // @[package.scala 32:76]
  assign _T_903_rs2 = _T_902 ? io_in[24:20] : _T_901_rs2; // @[package.scala 32:76]
  assign _T_903_rs3 = _T_902 ? io_in[31:27] : _T_901_rs3; // @[package.scala 32:76]
  assign _T_904 = _T_843 == 5'h1f; // @[package.scala 32:86]
  assign io_out_bits = _T_904 ? io_in : _T_903_bits; // @[RVC.scala 165:12]
  assign io_out_rd = _T_904 ? io_in[11:7] : _T_903_rd; // @[RVC.scala 165:12]
  assign io_out_rs1 = _T_904 ? io_in[19:15] : _T_903_rs1; // @[RVC.scala 165:12]
  assign io_out_rs2 = _T_904 ? io_in[24:20] : _T_903_rs2; // @[RVC.scala 165:12]
  assign io_out_rs3 = _T_904 ? io_in[31:27] : _T_903_rs3; // @[RVC.scala 165:12]
  assign io_rvc = io_in[1:0] != 2'h3; // @[RVC.scala 164:12]
  assign RVCExpander_covSum = 30'h0;
  assign io_covSum = RVCExpander_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNToRaw_preMul(
  input  [1:0]  io_op,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  output [23:0] io_mulAddA,
  output [23:0] io_mulAddB,
  output [47:0] io_mulAddC,
  output        io_toPostMul_isSigNaNAny,
  output        io_toPostMul_isNaNAOrB,
  output        io_toPostMul_isInfA,
  output        io_toPostMul_isZeroA,
  output        io_toPostMul_isInfB,
  output        io_toPostMul_isZeroB,
  output        io_toPostMul_signProd,
  output        io_toPostMul_isNaNC,
  output        io_toPostMul_isInfC,
  output        io_toPostMul_isZeroC,
  output [9:0]  io_toPostMul_sExpSum,
  output        io_toPostMul_doSubMags,
  output        io_toPostMul_CIsDominant,
  output [4:0]  io_toPostMul_CDom_CAlignDist,
  output [25:0] io_toPostMul_highAlignedSigC,
  output        io_toPostMul_bit0AlignedSigC,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawA_sig; // @[Cat.scala 29:58]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawB_sig; // @[Cat.scala 29:58]
  wire  rawC_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_36; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawC_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawC_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawC_sig; // @[Cat.scala 29:58]
  wire  _T_48; // @[MulAddRecFN.scala 98:30]
  wire  signProd; // @[MulAddRecFN.scala 98:42]
  wire [10:0] _T_50; // @[MulAddRecFN.scala 101:19]
  wire [10:0] sExpAlignedProd; // @[MulAddRecFN.scala 101:32]
  wire  _T_53; // @[MulAddRecFN.scala 103:30]
  wire  doSubMags; // @[MulAddRecFN.scala 103:42]
  wire [10:0] _GEN_0; // @[MulAddRecFN.scala 107:42]
  wire [10:0] sNatCAlignDist; // @[MulAddRecFN.scala 107:42]
  wire [9:0] posNatCAlignDist; // @[MulAddRecFN.scala 108:42]
  wire  _T_57; // @[MulAddRecFN.scala 109:35]
  wire  _T_58; // @[MulAddRecFN.scala 109:69]
  wire  isMinCAlign; // @[MulAddRecFN.scala 109:50]
  wire  _T_60; // @[MulAddRecFN.scala 111:60]
  wire  _T_61; // @[MulAddRecFN.scala 111:39]
  wire  CIsDominant; // @[MulAddRecFN.scala 111:23]
  wire  _T_62; // @[MulAddRecFN.scala 115:34]
  wire [6:0] _T_64; // @[MulAddRecFN.scala 115:16]
  wire [6:0] CAlignDist; // @[MulAddRecFN.scala 113:12]
  wire [24:0] _T_66; // @[MulAddRecFN.scala 121:16]
  wire [52:0] _T_68; // @[Bitwise.scala 72:12]
  wire [77:0] _T_70; // @[MulAddRecFN.scala 123:11]
  wire [77:0] mainAlignedSigC; // @[MulAddRecFN.scala 123:17]
  wire [26:0] _T_71; // @[MulAddRecFN.scala 125:30]
  wire  _T_74; // @[primitives.scala 121:54]
  wire  _T_76; // @[primitives.scala 121:54]
  wire  _T_78; // @[primitives.scala 121:54]
  wire  _T_80; // @[primitives.scala 121:54]
  wire  _T_82; // @[primitives.scala 121:54]
  wire  _T_84; // @[primitives.scala 121:54]
  wire  _T_86; // @[primitives.scala 124:57]
  wire [6:0] _T_92; // @[primitives.scala 125:20]
  wire [32:0] _T_94; // @[primitives.scala 77:58]
  wire [5:0] _T_110; // @[Cat.scala 29:58]
  wire [6:0] _GEN_1; // @[MulAddRecFN.scala 125:68]
  wire [6:0] _T_111; // @[MulAddRecFN.scala 125:68]
  wire  reduced4CExtra; // @[MulAddRecFN.scala 133:11]
  wire  _T_114; // @[MulAddRecFN.scala 137:39]
  wire  _T_116; // @[MulAddRecFN.scala 137:44]
  wire  _T_118; // @[MulAddRecFN.scala 138:39]
  wire  _T_119; // @[MulAddRecFN.scala 138:44]
  wire  _T_120; // @[MulAddRecFN.scala 136:16]
  wire [74:0] _T_121; // @[Cat.scala 29:58]
  wire [75:0] alignedSigC; // @[Cat.scala 29:58]
  wire  _T_125; // @[common.scala 81:46]
  wire  _T_128; // @[common.scala 81:46]
  wire  _T_129; // @[MulAddRecFN.scala 149:32]
  wire  _T_132; // @[common.scala 81:46]
  wire [10:0] _T_137; // @[MulAddRecFN.scala 161:53]
  wire [10:0] _T_138; // @[MulAddRecFN.scala 161:12]
  wire [29:0] MulAddRecFNToRaw_preMul_covSum;
  assign rawA_isZero = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_isNaN = _T_4 & io_a[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_sExp = {1'b0,$signed(io_a[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_sig = {1'h0,~rawA_isZero,io_a[22:0]}; // @[Cat.scala 29:58]
  assign rawB_isZero = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_20 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_isNaN = _T_20 & io_b[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_sExp = {1'b0,$signed(io_b[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_sig = {1'h0,~rawB_isZero,io_b[22:0]}; // @[Cat.scala 29:58]
  assign rawC_isZero = io_c[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_36 = io_c[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawC_isNaN = _T_36 & io_c[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawC_sign = io_c[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawC_sExp = {1'b0,$signed(io_c[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawC_sig = {1'h0,~rawC_isZero,io_c[22:0]}; // @[Cat.scala 29:58]
  assign _T_48 = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30]
  assign signProd = _T_48 ^ io_op[1]; // @[MulAddRecFN.scala 98:42]
  assign _T_50 = $signed(rawA_sExp) + $signed(rawB_sExp); // @[MulAddRecFN.scala 101:19]
  assign sExpAlignedProd = $signed(_T_50) + -11'she5; // @[MulAddRecFN.scala 101:32]
  assign _T_53 = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30]
  assign doSubMags = _T_53 ^ io_op[0]; // @[MulAddRecFN.scala 103:42]
  assign _GEN_0 = {{1{rawC_sExp[9]}},rawC_sExp}; // @[MulAddRecFN.scala 107:42]
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42]
  assign posNatCAlignDist = sNatCAlignDist[9:0]; // @[MulAddRecFN.scala 108:42]
  assign _T_57 = rawA_isZero | rawB_isZero; // @[MulAddRecFN.scala 109:35]
  assign _T_58 = $signed(sNatCAlignDist) < 11'sh0; // @[MulAddRecFN.scala 109:69]
  assign isMinCAlign = _T_57 | _T_58; // @[MulAddRecFN.scala 109:50]
  assign _T_60 = posNatCAlignDist <= 10'h18; // @[MulAddRecFN.scala 111:60]
  assign _T_61 = isMinCAlign | _T_60; // @[MulAddRecFN.scala 111:39]
  assign CIsDominant = ~rawC_isZero & _T_61; // @[MulAddRecFN.scala 111:23]
  assign _T_62 = posNatCAlignDist < 10'h4a; // @[MulAddRecFN.scala 115:34]
  assign _T_64 = _T_62 ? posNatCAlignDist[6:0] : 7'h4a; // @[MulAddRecFN.scala 115:16]
  assign CAlignDist = isMinCAlign ? 7'h0 : _T_64; // @[MulAddRecFN.scala 113:12]
  assign _T_66 = doSubMags ? ~rawC_sig : rawC_sig; // @[MulAddRecFN.scala 121:16]
  assign _T_68 = doSubMags ? 53'h1fffffffffffff : 53'h0; // @[Bitwise.scala 72:12]
  assign _T_70 = {_T_66,_T_68}; // @[MulAddRecFN.scala 123:11]
  assign mainAlignedSigC = $signed(_T_70) >>> CAlignDist; // @[MulAddRecFN.scala 123:17]
  assign _T_71 = {rawC_sig, 2'h0}; // @[MulAddRecFN.scala 125:30]
  assign _T_74 = |_T_71[3:0]; // @[primitives.scala 121:54]
  assign _T_76 = |_T_71[7:4]; // @[primitives.scala 121:54]
  assign _T_78 = |_T_71[11:8]; // @[primitives.scala 121:54]
  assign _T_80 = |_T_71[15:12]; // @[primitives.scala 121:54]
  assign _T_82 = |_T_71[19:16]; // @[primitives.scala 121:54]
  assign _T_84 = |_T_71[23:20]; // @[primitives.scala 121:54]
  assign _T_86 = |_T_71[26:24]; // @[primitives.scala 124:57]
  assign _T_92 = {_T_86,_T_84,_T_82,_T_80,_T_78,_T_76,_T_74}; // @[primitives.scala 125:20]
  assign _T_94 = -33'sh100000000 >>> CAlignDist[6:2]; // @[primitives.scala 77:58]
  assign _T_110 = {_T_94[14],_T_94[15],_T_94[16],_T_94[17],_T_94[18],_T_94[19]}; // @[Cat.scala 29:58]
  assign _GEN_1 = {{1'd0}, _T_110}; // @[MulAddRecFN.scala 125:68]
  assign _T_111 = _T_92 & _GEN_1; // @[MulAddRecFN.scala 125:68]
  assign reduced4CExtra = |_T_111; // @[MulAddRecFN.scala 133:11]
  assign _T_114 = &mainAlignedSigC[2:0]; // @[MulAddRecFN.scala 137:39]
  assign _T_116 = _T_114 & ~reduced4CExtra; // @[MulAddRecFN.scala 137:44]
  assign _T_118 = |mainAlignedSigC[2:0]; // @[MulAddRecFN.scala 138:39]
  assign _T_119 = _T_118 | reduced4CExtra; // @[MulAddRecFN.scala 138:44]
  assign _T_120 = doSubMags ? _T_116 : _T_119; // @[MulAddRecFN.scala 136:16]
  assign _T_121 = mainAlignedSigC[77:3]; // @[Cat.scala 29:58]
  assign alignedSigC = {_T_121,_T_120}; // @[Cat.scala 29:58]
  assign _T_125 = rawA_isNaN & ~rawA_sig[22]; // @[common.scala 81:46]
  assign _T_128 = rawB_isNaN & ~rawB_sig[22]; // @[common.scala 81:46]
  assign _T_129 = _T_125 | _T_128; // @[MulAddRecFN.scala 149:32]
  assign _T_132 = rawC_isNaN & ~rawC_sig[22]; // @[common.scala 81:46]
  assign _T_137 = $signed(sExpAlignedProd) - 11'sh18; // @[MulAddRecFN.scala 161:53]
  assign _T_138 = CIsDominant ? $signed({{1{rawC_sExp[9]}},rawC_sExp}) : $signed(_T_137); // @[MulAddRecFN.scala 161:12]
  assign io_mulAddA = rawA_sig[23:0]; // @[MulAddRecFN.scala 144:16]
  assign io_mulAddB = rawB_sig[23:0]; // @[MulAddRecFN.scala 145:16]
  assign io_mulAddC = alignedSigC[48:1]; // @[MulAddRecFN.scala 146:16]
  assign io_toPostMul_isSigNaNAny = _T_129 | _T_132; // @[MulAddRecFN.scala 148:30]
  assign io_toPostMul_isNaNAOrB = rawA_isNaN | rawB_isNaN; // @[MulAddRecFN.scala 151:28]
  assign io_toPostMul_isInfA = _T_4 & ~io_a[29]; // @[MulAddRecFN.scala 152:28]
  assign io_toPostMul_isZeroA = io_a[31:29] == 3'h0; // @[MulAddRecFN.scala 153:28]
  assign io_toPostMul_isInfB = _T_20 & ~io_b[29]; // @[MulAddRecFN.scala 154:28]
  assign io_toPostMul_isZeroB = io_b[31:29] == 3'h0; // @[MulAddRecFN.scala 155:28]
  assign io_toPostMul_signProd = _T_48 ^ io_op[1]; // @[MulAddRecFN.scala 156:28]
  assign io_toPostMul_isNaNC = _T_36 & io_c[29]; // @[MulAddRecFN.scala 157:28]
  assign io_toPostMul_isInfC = _T_36 & ~io_c[29]; // @[MulAddRecFN.scala 158:28]
  assign io_toPostMul_isZeroC = io_c[31:29] == 3'h0; // @[MulAddRecFN.scala 159:28]
  assign io_toPostMul_sExpSum = _T_138[9:0]; // @[MulAddRecFN.scala 160:28]
  assign io_toPostMul_doSubMags = _T_53 ^ io_op[0]; // @[MulAddRecFN.scala 162:28]
  assign io_toPostMul_CIsDominant = ~rawC_isZero & _T_61; // @[MulAddRecFN.scala 163:30]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[4:0]; // @[MulAddRecFN.scala 164:34]
  assign io_toPostMul_highAlignedSigC = alignedSigC[74:49]; // @[MulAddRecFN.scala 165:34]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:34]
  assign MulAddRecFNToRaw_preMul_covSum = 30'h0;
  assign io_covSum = MulAddRecFNToRaw_preMul_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNToRaw_postMul(
  input         io_fromPreMul_isSigNaNAny,
  input         io_fromPreMul_isNaNAOrB,
  input         io_fromPreMul_isInfA,
  input         io_fromPreMul_isZeroA,
  input         io_fromPreMul_isInfB,
  input         io_fromPreMul_isZeroB,
  input         io_fromPreMul_signProd,
  input         io_fromPreMul_isNaNC,
  input         io_fromPreMul_isInfC,
  input         io_fromPreMul_isZeroC,
  input  [9:0]  io_fromPreMul_sExpSum,
  input         io_fromPreMul_doSubMags,
  input         io_fromPreMul_CIsDominant,
  input  [4:0]  io_fromPreMul_CDom_CAlignDist,
  input  [25:0] io_fromPreMul_highAlignedSigC,
  input         io_fromPreMul_bit0AlignedSigC,
  input  [48:0] io_mulAddResult,
  input  [2:0]  io_roundingMode,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_min; // @[MulAddRecFN.scala 188:45]
  wire  CDom_sign; // @[MulAddRecFN.scala 192:42]
  wire [25:0] _T_2; // @[MulAddRecFN.scala 195:47]
  wire [25:0] _T_3; // @[MulAddRecFN.scala 194:16]
  wire [74:0] sigSum; // @[Cat.scala 29:58]
  wire [1:0] _T_6; // @[MulAddRecFN.scala 205:69]
  wire [9:0] _GEN_0; // @[MulAddRecFN.scala 205:43]
  wire [9:0] CDom_sExp; // @[MulAddRecFN.scala 205:43]
  wire [49:0] _T_14; // @[Cat.scala 29:58]
  wire [49:0] CDom_absSigSum; // @[MulAddRecFN.scala 207:12]
  wire  _T_17; // @[MulAddRecFN.scala 217:36]
  wire  _T_19; // @[MulAddRecFN.scala 218:37]
  wire  CDom_absSigSumExtra; // @[MulAddRecFN.scala 216:12]
  wire [80:0] _GEN_1; // @[MulAddRecFN.scala 221:24]
  wire [80:0] _T_20; // @[MulAddRecFN.scala 221:24]
  wire [28:0] CDom_mainSig; // @[MulAddRecFN.scala 221:56]
  wire [26:0] _T_22; // @[MulAddRecFN.scala 224:53]
  wire  _T_25; // @[primitives.scala 121:54]
  wire  _T_27; // @[primitives.scala 121:54]
  wire  _T_29; // @[primitives.scala 121:54]
  wire  _T_31; // @[primitives.scala 121:54]
  wire  _T_33; // @[primitives.scala 121:54]
  wire  _T_35; // @[primitives.scala 121:54]
  wire  _T_37; // @[primitives.scala 124:57]
  wire [6:0] _T_43; // @[primitives.scala 125:20]
  wire [8:0] _T_46; // @[primitives.scala 77:58]
  wire [5:0] _T_62; // @[Cat.scala 29:58]
  wire [6:0] _GEN_2; // @[MulAddRecFN.scala 224:72]
  wire [6:0] _T_63; // @[MulAddRecFN.scala 224:72]
  wire  CDom_reduced4SigExtra; // @[MulAddRecFN.scala 225:73]
  wire  _T_66; // @[MulAddRecFN.scala 228:32]
  wire  _T_67; // @[MulAddRecFN.scala 228:36]
  wire  _T_68; // @[MulAddRecFN.scala 228:61]
  wire [26:0] CDom_sig; // @[Cat.scala 29:58]
  wire  notCDom_signSigSum; // @[MulAddRecFN.scala 234:36]
  wire [50:0] _GEN_3; // @[MulAddRecFN.scala 238:41]
  wire [50:0] _T_73; // @[MulAddRecFN.scala 238:41]
  wire [50:0] notCDom_absSigSum; // @[MulAddRecFN.scala 236:12]
  wire  _T_76; // @[primitives.scala 104:54]
  wire  _T_78; // @[primitives.scala 104:54]
  wire  _T_80; // @[primitives.scala 104:54]
  wire  _T_82; // @[primitives.scala 104:54]
  wire  _T_84; // @[primitives.scala 104:54]
  wire  _T_86; // @[primitives.scala 104:54]
  wire  _T_88; // @[primitives.scala 104:54]
  wire  _T_90; // @[primitives.scala 104:54]
  wire  _T_92; // @[primitives.scala 104:54]
  wire  _T_94; // @[primitives.scala 104:54]
  wire  _T_96; // @[primitives.scala 104:54]
  wire  _T_98; // @[primitives.scala 104:54]
  wire  _T_100; // @[primitives.scala 104:54]
  wire  _T_102; // @[primitives.scala 104:54]
  wire  _T_104; // @[primitives.scala 104:54]
  wire  _T_106; // @[primitives.scala 104:54]
  wire  _T_108; // @[primitives.scala 104:54]
  wire  _T_110; // @[primitives.scala 104:54]
  wire  _T_112; // @[primitives.scala 104:54]
  wire  _T_114; // @[primitives.scala 104:54]
  wire  _T_116; // @[primitives.scala 104:54]
  wire  _T_118; // @[primitives.scala 104:54]
  wire  _T_120; // @[primitives.scala 104:54]
  wire  _T_122; // @[primitives.scala 104:54]
  wire  _T_124; // @[primitives.scala 104:54]
  wire  _T_126; // @[primitives.scala 107:57]
  wire [5:0] _T_131; // @[primitives.scala 108:20]
  wire [12:0] _T_138; // @[primitives.scala 108:20]
  wire [5:0] _T_143; // @[primitives.scala 108:20]
  wire [25:0] notCDom_reduced2AbsSigSum; // @[primitives.scala 108:20]
  wire [4:0] _T_177; // @[Mux.scala 47:69]
  wire [4:0] _T_178; // @[Mux.scala 47:69]
  wire [4:0] _T_179; // @[Mux.scala 47:69]
  wire [4:0] _T_180; // @[Mux.scala 47:69]
  wire [4:0] _T_181; // @[Mux.scala 47:69]
  wire [4:0] _T_182; // @[Mux.scala 47:69]
  wire [4:0] _T_183; // @[Mux.scala 47:69]
  wire [4:0] _T_184; // @[Mux.scala 47:69]
  wire [4:0] _T_185; // @[Mux.scala 47:69]
  wire [4:0] _T_186; // @[Mux.scala 47:69]
  wire [4:0] _T_187; // @[Mux.scala 47:69]
  wire [4:0] _T_188; // @[Mux.scala 47:69]
  wire [4:0] _T_189; // @[Mux.scala 47:69]
  wire [4:0] _T_190; // @[Mux.scala 47:69]
  wire [4:0] _T_191; // @[Mux.scala 47:69]
  wire [4:0] _T_192; // @[Mux.scala 47:69]
  wire [4:0] _T_193; // @[Mux.scala 47:69]
  wire [4:0] _T_194; // @[Mux.scala 47:69]
  wire [4:0] _T_195; // @[Mux.scala 47:69]
  wire [4:0] _T_196; // @[Mux.scala 47:69]
  wire [4:0] _T_197; // @[Mux.scala 47:69]
  wire [4:0] _T_198; // @[Mux.scala 47:69]
  wire [4:0] _T_199; // @[Mux.scala 47:69]
  wire [4:0] _T_200; // @[Mux.scala 47:69]
  wire [4:0] notCDom_normDistReduced2; // @[Mux.scala 47:69]
  wire [5:0] notCDom_nearNormDist; // @[MulAddRecFN.scala 242:56]
  wire [6:0] _T_201; // @[MulAddRecFN.scala 243:69]
  wire [9:0] _GEN_4; // @[MulAddRecFN.scala 243:46]
  wire [9:0] notCDom_sExp; // @[MulAddRecFN.scala 243:46]
  wire [113:0] _GEN_5; // @[MulAddRecFN.scala 245:27]
  wire [113:0] _T_204; // @[MulAddRecFN.scala 245:27]
  wire [28:0] notCDom_mainSig; // @[MulAddRecFN.scala 245:50]
  wire  _T_209; // @[primitives.scala 104:54]
  wire  _T_211; // @[primitives.scala 104:54]
  wire  _T_213; // @[primitives.scala 104:54]
  wire  _T_215; // @[primitives.scala 104:54]
  wire  _T_217; // @[primitives.scala 104:54]
  wire  _T_219; // @[primitives.scala 104:54]
  wire  _T_221; // @[primitives.scala 107:57]
  wire [6:0] _T_227; // @[primitives.scala 108:20]
  wire [16:0] _T_230; // @[primitives.scala 77:58]
  wire [5:0] _T_246; // @[Cat.scala 29:58]
  wire [6:0] _GEN_6; // @[MulAddRecFN.scala 249:78]
  wire [6:0] _T_247; // @[MulAddRecFN.scala 249:78]
  wire  notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 251:11]
  wire  _T_250; // @[MulAddRecFN.scala 254:35]
  wire  _T_251; // @[MulAddRecFN.scala 254:39]
  wire [26:0] notCDom_sig; // @[Cat.scala 29:58]
  wire  notCDom_completeCancellation; // @[MulAddRecFN.scala 257:50]
  wire  _T_253; // @[MulAddRecFN.scala 261:36]
  wire  notCDom_sign; // @[MulAddRecFN.scala 259:12]
  wire  notNaN_isInfProd; // @[MulAddRecFN.scala 266:49]
  wire  notNaN_isInfOut; // @[MulAddRecFN.scala 267:44]
  wire  _T_254; // @[MulAddRecFN.scala 269:32]
  wire  notNaN_addZeros; // @[MulAddRecFN.scala 269:58]
  wire  _T_255; // @[MulAddRecFN.scala 274:31]
  wire  _T_256; // @[MulAddRecFN.scala 273:35]
  wire  _T_257; // @[MulAddRecFN.scala 275:32]
  wire  _T_258; // @[MulAddRecFN.scala 274:57]
  wire  _T_261; // @[MulAddRecFN.scala 276:36]
  wire  _T_262; // @[MulAddRecFN.scala 277:61]
  wire  _T_263; // @[MulAddRecFN.scala 278:35]
  wire  _T_267; // @[MulAddRecFN.scala 285:42]
  wire  _T_269; // @[MulAddRecFN.scala 287:27]
  wire  _T_270; // @[MulAddRecFN.scala 288:31]
  wire  _T_271; // @[MulAddRecFN.scala 287:54]
  wire  _T_273; // @[MulAddRecFN.scala 289:26]
  wire  _T_274; // @[MulAddRecFN.scala 289:48]
  wire  _T_275; // @[MulAddRecFN.scala 290:36]
  wire  _T_276; // @[MulAddRecFN.scala 288:43]
  wire  _T_277; // @[MulAddRecFN.scala 291:26]
  wire  _T_278; // @[MulAddRecFN.scala 292:37]
  wire  _T_279; // @[MulAddRecFN.scala 291:46]
  wire  _T_280; // @[MulAddRecFN.scala 290:48]
  wire  _T_283; // @[MulAddRecFN.scala 293:28]
  wire  _T_284; // @[MulAddRecFN.scala 294:17]
  wire  _T_285; // @[MulAddRecFN.scala 293:49]
  wire [29:0] MulAddRecFNToRaw_postMul_covSum;
  assign roundingMode_min = io_roundingMode == 3'h2; // @[MulAddRecFN.scala 188:45]
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42]
  assign _T_2 = io_fromPreMul_highAlignedSigC + 26'h1; // @[MulAddRecFN.scala 195:47]
  assign _T_3 = io_mulAddResult[48] ? _T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16]
  assign sigSum = {_T_3,io_mulAddResult[47:0],io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 29:58]
  assign _T_6 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69]
  assign _GEN_0 = {{8{_T_6[1]}},_T_6}; // @[MulAddRecFN.scala 205:43]
  assign CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43]
  assign _T_14 = {1'h0,io_fromPreMul_highAlignedSigC[25:24],sigSum[72:26]}; // @[Cat.scala 29:58]
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? ~sigSum[74:25] : _T_14; // @[MulAddRecFN.scala 207:12]
  assign _T_17 = |~sigSum[24:1]; // @[MulAddRecFN.scala 217:36]
  assign _T_19 = |sigSum[25:1]; // @[MulAddRecFN.scala 218:37]
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_17 : _T_19; // @[MulAddRecFN.scala 216:12]
  assign _GEN_1 = {{31'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24]
  assign _T_20 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24]
  assign CDom_mainSig = _T_20[49:21]; // @[MulAddRecFN.scala 221:56]
  assign _T_22 = {CDom_absSigSum[23:0], 3'h0}; // @[MulAddRecFN.scala 224:53]
  assign _T_25 = |_T_22[3:0]; // @[primitives.scala 121:54]
  assign _T_27 = |_T_22[7:4]; // @[primitives.scala 121:54]
  assign _T_29 = |_T_22[11:8]; // @[primitives.scala 121:54]
  assign _T_31 = |_T_22[15:12]; // @[primitives.scala 121:54]
  assign _T_33 = |_T_22[19:16]; // @[primitives.scala 121:54]
  assign _T_35 = |_T_22[23:20]; // @[primitives.scala 121:54]
  assign _T_37 = |_T_22[26:24]; // @[primitives.scala 124:57]
  assign _T_43 = {_T_37,_T_35,_T_33,_T_31,_T_29,_T_27,_T_25}; // @[primitives.scala 125:20]
  assign _T_46 = -9'sh100 >>> ~io_fromPreMul_CDom_CAlignDist[4:2]; // @[primitives.scala 77:58]
  assign _T_62 = {_T_46[1],_T_46[2],_T_46[3],_T_46[4],_T_46[5],_T_46[6]}; // @[Cat.scala 29:58]
  assign _GEN_2 = {{1'd0}, _T_62}; // @[MulAddRecFN.scala 224:72]
  assign _T_63 = _T_43 & _GEN_2; // @[MulAddRecFN.scala 224:72]
  assign CDom_reduced4SigExtra = |_T_63; // @[MulAddRecFN.scala 225:73]
  assign _T_66 = |CDom_mainSig[2:0]; // @[MulAddRecFN.scala 228:32]
  assign _T_67 = _T_66 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36]
  assign _T_68 = _T_67 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61]
  assign CDom_sig = {CDom_mainSig[28:3],_T_68}; // @[Cat.scala 29:58]
  assign notCDom_signSigSum = sigSum[51]; // @[MulAddRecFN.scala 234:36]
  assign _GEN_3 = {{50'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41]
  assign _T_73 = sigSum[50:0] + _GEN_3; // @[MulAddRecFN.scala 238:41]
  assign notCDom_absSigSum = notCDom_signSigSum ? ~sigSum[50:0] : _T_73; // @[MulAddRecFN.scala 236:12]
  assign _T_76 = |notCDom_absSigSum[1:0]; // @[primitives.scala 104:54]
  assign _T_78 = |notCDom_absSigSum[3:2]; // @[primitives.scala 104:54]
  assign _T_80 = |notCDom_absSigSum[5:4]; // @[primitives.scala 104:54]
  assign _T_82 = |notCDom_absSigSum[7:6]; // @[primitives.scala 104:54]
  assign _T_84 = |notCDom_absSigSum[9:8]; // @[primitives.scala 104:54]
  assign _T_86 = |notCDom_absSigSum[11:10]; // @[primitives.scala 104:54]
  assign _T_88 = |notCDom_absSigSum[13:12]; // @[primitives.scala 104:54]
  assign _T_90 = |notCDom_absSigSum[15:14]; // @[primitives.scala 104:54]
  assign _T_92 = |notCDom_absSigSum[17:16]; // @[primitives.scala 104:54]
  assign _T_94 = |notCDom_absSigSum[19:18]; // @[primitives.scala 104:54]
  assign _T_96 = |notCDom_absSigSum[21:20]; // @[primitives.scala 104:54]
  assign _T_98 = |notCDom_absSigSum[23:22]; // @[primitives.scala 104:54]
  assign _T_100 = |notCDom_absSigSum[25:24]; // @[primitives.scala 104:54]
  assign _T_102 = |notCDom_absSigSum[27:26]; // @[primitives.scala 104:54]
  assign _T_104 = |notCDom_absSigSum[29:28]; // @[primitives.scala 104:54]
  assign _T_106 = |notCDom_absSigSum[31:30]; // @[primitives.scala 104:54]
  assign _T_108 = |notCDom_absSigSum[33:32]; // @[primitives.scala 104:54]
  assign _T_110 = |notCDom_absSigSum[35:34]; // @[primitives.scala 104:54]
  assign _T_112 = |notCDom_absSigSum[37:36]; // @[primitives.scala 104:54]
  assign _T_114 = |notCDom_absSigSum[39:38]; // @[primitives.scala 104:54]
  assign _T_116 = |notCDom_absSigSum[41:40]; // @[primitives.scala 104:54]
  assign _T_118 = |notCDom_absSigSum[43:42]; // @[primitives.scala 104:54]
  assign _T_120 = |notCDom_absSigSum[45:44]; // @[primitives.scala 104:54]
  assign _T_122 = |notCDom_absSigSum[47:46]; // @[primitives.scala 104:54]
  assign _T_124 = |notCDom_absSigSum[49:48]; // @[primitives.scala 104:54]
  assign _T_126 = |notCDom_absSigSum[50]; // @[primitives.scala 107:57]
  assign _T_131 = {_T_86,_T_84,_T_82,_T_80,_T_78,_T_76}; // @[primitives.scala 108:20]
  assign _T_138 = {_T_100,_T_98,_T_96,_T_94,_T_92,_T_90,_T_88,_T_131}; // @[primitives.scala 108:20]
  assign _T_143 = {_T_112,_T_110,_T_108,_T_106,_T_104,_T_102}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum = {_T_126,_T_124,_T_122,_T_120,_T_118,_T_116,_T_114,_T_143,_T_138}; // @[primitives.scala 108:20]
  assign _T_177 = notCDom_reduced2AbsSigSum[1] ? 5'h18 : 5'h19; // @[Mux.scala 47:69]
  assign _T_178 = notCDom_reduced2AbsSigSum[2] ? 5'h17 : _T_177; // @[Mux.scala 47:69]
  assign _T_179 = notCDom_reduced2AbsSigSum[3] ? 5'h16 : _T_178; // @[Mux.scala 47:69]
  assign _T_180 = notCDom_reduced2AbsSigSum[4] ? 5'h15 : _T_179; // @[Mux.scala 47:69]
  assign _T_181 = notCDom_reduced2AbsSigSum[5] ? 5'h14 : _T_180; // @[Mux.scala 47:69]
  assign _T_182 = notCDom_reduced2AbsSigSum[6] ? 5'h13 : _T_181; // @[Mux.scala 47:69]
  assign _T_183 = notCDom_reduced2AbsSigSum[7] ? 5'h12 : _T_182; // @[Mux.scala 47:69]
  assign _T_184 = notCDom_reduced2AbsSigSum[8] ? 5'h11 : _T_183; // @[Mux.scala 47:69]
  assign _T_185 = notCDom_reduced2AbsSigSum[9] ? 5'h10 : _T_184; // @[Mux.scala 47:69]
  assign _T_186 = notCDom_reduced2AbsSigSum[10] ? 5'hf : _T_185; // @[Mux.scala 47:69]
  assign _T_187 = notCDom_reduced2AbsSigSum[11] ? 5'he : _T_186; // @[Mux.scala 47:69]
  assign _T_188 = notCDom_reduced2AbsSigSum[12] ? 5'hd : _T_187; // @[Mux.scala 47:69]
  assign _T_189 = notCDom_reduced2AbsSigSum[13] ? 5'hc : _T_188; // @[Mux.scala 47:69]
  assign _T_190 = notCDom_reduced2AbsSigSum[14] ? 5'hb : _T_189; // @[Mux.scala 47:69]
  assign _T_191 = notCDom_reduced2AbsSigSum[15] ? 5'ha : _T_190; // @[Mux.scala 47:69]
  assign _T_192 = notCDom_reduced2AbsSigSum[16] ? 5'h9 : _T_191; // @[Mux.scala 47:69]
  assign _T_193 = notCDom_reduced2AbsSigSum[17] ? 5'h8 : _T_192; // @[Mux.scala 47:69]
  assign _T_194 = notCDom_reduced2AbsSigSum[18] ? 5'h7 : _T_193; // @[Mux.scala 47:69]
  assign _T_195 = notCDom_reduced2AbsSigSum[19] ? 5'h6 : _T_194; // @[Mux.scala 47:69]
  assign _T_196 = notCDom_reduced2AbsSigSum[20] ? 5'h5 : _T_195; // @[Mux.scala 47:69]
  assign _T_197 = notCDom_reduced2AbsSigSum[21] ? 5'h4 : _T_196; // @[Mux.scala 47:69]
  assign _T_198 = notCDom_reduced2AbsSigSum[22] ? 5'h3 : _T_197; // @[Mux.scala 47:69]
  assign _T_199 = notCDom_reduced2AbsSigSum[23] ? 5'h2 : _T_198; // @[Mux.scala 47:69]
  assign _T_200 = notCDom_reduced2AbsSigSum[24] ? 5'h1 : _T_199; // @[Mux.scala 47:69]
  assign notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[25] ? 5'h0 : _T_200; // @[Mux.scala 47:69]
  assign notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56]
  assign _T_201 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69]
  assign _GEN_4 = {{3{_T_201[6]}},_T_201}; // @[MulAddRecFN.scala 243:46]
  assign notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_4); // @[MulAddRecFN.scala 243:46]
  assign _GEN_5 = {{63'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27]
  assign _T_204 = _GEN_5 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27]
  assign notCDom_mainSig = _T_204[51:23]; // @[MulAddRecFN.scala 245:50]
  assign _T_209 = |notCDom_reduced2AbsSigSum[1:0]; // @[primitives.scala 104:54]
  assign _T_211 = |notCDom_reduced2AbsSigSum[3:2]; // @[primitives.scala 104:54]
  assign _T_213 = |notCDom_reduced2AbsSigSum[5:4]; // @[primitives.scala 104:54]
  assign _T_215 = |notCDom_reduced2AbsSigSum[7:6]; // @[primitives.scala 104:54]
  assign _T_217 = |notCDom_reduced2AbsSigSum[9:8]; // @[primitives.scala 104:54]
  assign _T_219 = |notCDom_reduced2AbsSigSum[11:10]; // @[primitives.scala 104:54]
  assign _T_221 = |notCDom_reduced2AbsSigSum[12]; // @[primitives.scala 107:57]
  assign _T_227 = {_T_221,_T_219,_T_217,_T_215,_T_213,_T_211,_T_209}; // @[primitives.scala 108:20]
  assign _T_230 = -17'sh10000 >>> ~notCDom_normDistReduced2[4:1]; // @[primitives.scala 77:58]
  assign _T_246 = {_T_230[1],_T_230[2],_T_230[3],_T_230[4],_T_230[5],_T_230[6]}; // @[Cat.scala 29:58]
  assign _GEN_6 = {{1'd0}, _T_246}; // @[MulAddRecFN.scala 249:78]
  assign _T_247 = _T_227 & _GEN_6; // @[MulAddRecFN.scala 249:78]
  assign notCDom_reduced4SigExtra = |_T_247; // @[MulAddRecFN.scala 251:11]
  assign _T_250 = |notCDom_mainSig[2:0]; // @[MulAddRecFN.scala 254:35]
  assign _T_251 = _T_250 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39]
  assign notCDom_sig = {notCDom_mainSig[28:3],_T_251}; // @[Cat.scala 29:58]
  assign notCDom_completeCancellation = notCDom_sig[26:25] == 2'h0; // @[MulAddRecFN.scala 257:50]
  assign _T_253 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36]
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _T_253; // @[MulAddRecFN.scala 259:12]
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49]
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  assign _T_254 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32]
  assign notNaN_addZeros = _T_254 & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58]
  assign _T_255 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31]
  assign _T_256 = io_fromPreMul_isSigNaNAny | _T_255; // @[MulAddRecFN.scala 273:35]
  assign _T_257 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32]
  assign _T_258 = _T_256 | _T_257; // @[MulAddRecFN.scala 274:57]
  assign _T_261 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36]
  assign _T_262 = _T_261 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61]
  assign _T_263 = _T_262 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35]
  assign _T_267 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42]
  assign _T_269 = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27]
  assign _T_270 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31]
  assign _T_271 = _T_269 | _T_270; // @[MulAddRecFN.scala 287:54]
  assign _T_273 = notNaN_addZeros & ~roundingMode_min; // @[MulAddRecFN.scala 289:26]
  assign _T_274 = _T_273 & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48]
  assign _T_275 = _T_274 & CDom_sign; // @[MulAddRecFN.scala 290:36]
  assign _T_276 = _T_271 | _T_275; // @[MulAddRecFN.scala 288:43]
  assign _T_277 = notNaN_addZeros & roundingMode_min; // @[MulAddRecFN.scala 291:26]
  assign _T_278 = io_fromPreMul_signProd | CDom_sign; // @[MulAddRecFN.scala 292:37]
  assign _T_279 = _T_277 & _T_278; // @[MulAddRecFN.scala 291:46]
  assign _T_280 = _T_276 | _T_279; // @[MulAddRecFN.scala 290:48]
  assign _T_283 = ~notNaN_isInfOut & ~notNaN_addZeros; // @[MulAddRecFN.scala 293:28]
  assign _T_284 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17]
  assign _T_285 = _T_283 & _T_284; // @[MulAddRecFN.scala 293:49]
  assign io_invalidExc = _T_258 | _T_263; // @[MulAddRecFN.scala 272:19]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21]
  assign io_rawOut_isZero = notNaN_addZeros | _T_267; // @[MulAddRecFN.scala 283:22]
  assign io_rawOut_sign = _T_280 | _T_285; // @[MulAddRecFN.scala 286:20]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19]
  assign MulAddRecFNToRaw_postMul_covSum = 30'h0;
  assign io_covSum = MulAddRecFNToRaw_postMul_covSum;
  assign metaAssert = 1'h0;
endmodule
module RoundAnyRawFNToRecFN_1(
  input         io_in_isZero,
  input         io_in_sign,
  input  [8:0]  io_in_sExp,
  input  [64:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire [9:0] _T_3; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [9:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 104:31]
  wire  _T_7; // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [26:0] adjustedSig; // @[Cat.scala 29:58]
  wire [26:0] _T_14; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_15; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _T_16; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_17; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_19; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_20; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_21; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_22; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [26:0] _T_23; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _T_25; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_26; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_28; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [25:0] _T_30; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _T_32; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _T_34; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_36; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [25:0] _T_38; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [25:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_39; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_40; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_42; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [9:0] _GEN_1; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [10:0] _T_43; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:64]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire [8:0] _T_75; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [9:0] _T_101; // @[Cat.scala 29:58]
  wire [1:0] _T_103; // @[Cat.scala 29:58]
  wire [29:0] RoundAnyRawFNToRecFN_1_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign _T_3 = $signed(io_in_sExp) + 9'sh80; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign sAdjustedExp = {1'b0,$signed(_T_3[8:0])}; // @[RoundAnyRawFNToRecFN.scala 104:31]
  assign _T_7 = |io_in_sig[38:0]; // @[RoundAnyRawFNToRecFN.scala 115:60]
  assign adjustedSig = {io_in_sig[64:39],_T_7}; // @[Cat.scala 29:58]
  assign _T_14 = adjustedSig & 27'h2; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_15 = |_T_14; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_16 = adjustedSig & 27'h1; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_17 = |_T_16; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign common_inexact = _T_15 | _T_17; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_19 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_20 = _T_19 & _T_15; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_21 = roundMagUp & common_inexact; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_22 = _T_20 | _T_21; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_23 = adjustedSig | 27'h3; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_25 = _T_23[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_26 = roundingMode_near_even & _T_15; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_28 = _T_26 & ~_T_17; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_30 = _T_28 ? 26'h1 : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_32 = _T_25 & ~_T_30; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_34 = adjustedSig & 27'h7fffffc; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_36 = roundingMode_odd & common_inexact; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_38 = _T_36 ? 26'h1 : 26'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_0 = {{1'd0}, _T_34[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_39 = _GEN_0 | _T_38; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_40 = _T_22 ? _T_32 : _T_39; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_42 = {1'b0,$signed(_T_40[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_1 = {{7{_T_42[2]}},_T_42}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_43 = $signed(sAdjustedExp) + $signed(_GEN_1); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_43[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = _T_40[22:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  assign commonCase = ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:64]
  assign inexact = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign _T_75 = io_in_isZero ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign expOut = common_expOut & ~_T_75; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign fractOut = io_in_isZero ? 23'h0 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_101 = {io_in_sign,expOut}; // @[Cat.scala 29:58]
  assign _T_103 = {1'h0,inexact}; // @[Cat.scala 29:58]
  assign io_out = {_T_101,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {3'h0,_T_103}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_1_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module RoundAnyRawFNToRecFN_2(
  input         io_in_isZero,
  input         io_in_sign,
  input  [8:0]  io_in_sExp,
  input  [64:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire [11:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [12:0] _T_3; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [12:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 104:31]
  wire  _T_7; // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [55:0] adjustedSig; // @[Cat.scala 29:58]
  wire [55:0] _T_14; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_15; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [55:0] _T_16; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_17; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_19; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_20; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_21; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_22; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [55:0] _T_23; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [54:0] _T_25; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_26; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_28; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [54:0] _T_30; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [54:0] _T_32; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [55:0] _T_34; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_36; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [54:0] _T_38; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [54:0] _GEN_1; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _T_39; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _T_40; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_42; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [12:0] _GEN_2; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [13:0] _T_43; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [11:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [51:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:64]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire [11:0] _T_75; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [11:0] expOut; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [51:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [12:0] _T_101; // @[Cat.scala 29:58]
  wire [1:0] _T_103; // @[Cat.scala 29:58]
  wire [29:0] RoundAnyRawFNToRecFN_2_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign _GEN_0 = {{3{io_in_sExp[8]}},io_in_sExp}; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign _T_3 = $signed(_GEN_0) + 12'sh780; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign sAdjustedExp = {1'b0,$signed(_T_3[11:0])}; // @[RoundAnyRawFNToRecFN.scala 104:31]
  assign _T_7 = |io_in_sig[9:0]; // @[RoundAnyRawFNToRecFN.scala 115:60]
  assign adjustedSig = {io_in_sig[64:10],_T_7}; // @[Cat.scala 29:58]
  assign _T_14 = adjustedSig & 56'h2; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_15 = |_T_14; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_16 = adjustedSig & 56'h1; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_17 = |_T_16; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign common_inexact = _T_15 | _T_17; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_19 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_20 = _T_19 & _T_15; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_21 = roundMagUp & common_inexact; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_22 = _T_20 | _T_21; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_23 = adjustedSig | 56'h3; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_25 = _T_23[55:2] + 54'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_26 = roundingMode_near_even & _T_15; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_28 = _T_26 & ~_T_17; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_30 = _T_28 ? 55'h1 : 55'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_32 = _T_25 & ~_T_30; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_34 = adjustedSig & 56'hfffffffffffffc; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_36 = roundingMode_odd & common_inexact; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_38 = _T_36 ? 55'h1 : 55'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_1 = {{1'd0}, _T_34[55:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_39 = _GEN_1 | _T_38; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_40 = _T_22 ? _T_32 : _T_39; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_42 = {1'b0,$signed(_T_40[54:53])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_2 = {{10{_T_42[2]}},_T_42}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_43 = $signed(sAdjustedExp) + $signed(_GEN_2); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_43[11:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = _T_40[51:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  assign commonCase = ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:64]
  assign inexact = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign _T_75 = io_in_isZero ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign expOut = common_expOut & ~_T_75; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign fractOut = io_in_isZero ? 52'h0 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_101 = {io_in_sign,expOut}; // @[Cat.scala 29:58]
  assign _T_103 = {1'h0,inexact}; // @[Cat.scala 29:58]
  assign io_out = {_T_101,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {3'h0,_T_103}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_2_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_2_covSum;
  assign metaAssert = 1'h0;
endmodule
module RoundAnyRawFNToRecFN_3(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [53:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire [13:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 108:24]
  wire  _T_5; // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [26:0] adjustedSig; // @[Cat.scala 29:58]
  wire  _T_8; // @[primitives.scala 57:25]
  wire  _T_10; // @[primitives.scala 57:25]
  wire  _T_12; // @[primitives.scala 57:25]
  wire [5:0] _T_13; // @[primitives.scala 58:26]
  wire [64:0] _T_14; // @[primitives.scala 77:58]
  wire [15:0] _T_20; // @[Bitwise.scala 103:31]
  wire [15:0] _T_22; // @[Bitwise.scala 103:65]
  wire [15:0] _T_24; // @[Bitwise.scala 103:75]
  wire [15:0] _T_25; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_0; // @[Bitwise.scala 103:31]
  wire [15:0] _T_30; // @[Bitwise.scala 103:31]
  wire [15:0] _T_32; // @[Bitwise.scala 103:65]
  wire [15:0] _T_34; // @[Bitwise.scala 103:75]
  wire [15:0] _T_35; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [15:0] _T_40; // @[Bitwise.scala 103:31]
  wire [15:0] _T_42; // @[Bitwise.scala 103:65]
  wire [15:0] _T_44; // @[Bitwise.scala 103:75]
  wire [15:0] _T_45; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [15:0] _T_50; // @[Bitwise.scala 103:31]
  wire [15:0] _T_52; // @[Bitwise.scala 103:65]
  wire [15:0] _T_54; // @[Bitwise.scala 103:75]
  wire [15:0] _T_55; // @[Bitwise.scala 103:39]
  wire [21:0] _T_72; // @[Cat.scala 29:58]
  wire [21:0] _T_74; // @[primitives.scala 74:21]
  wire [24:0] _T_76; // @[Cat.scala 29:58]
  wire [2:0] _T_86; // @[Cat.scala 29:58]
  wire [2:0] _T_87; // @[primitives.scala 61:24]
  wire [24:0] _T_88; // @[primitives.scala 66:24]
  wire [24:0] _T_89; // @[primitives.scala 61:24]
  wire [26:0] _T_91; // @[Cat.scala 29:58]
  wire [26:0] _T_93; // @[Cat.scala 29:58]
  wire [26:0] _T_95; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [26:0] _T_96; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_97; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _T_98; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_99; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  _T_100; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_101; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_102; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_103; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_104; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [26:0] _T_105; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _T_107; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_108; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_110; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [25:0] _T_112; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _T_114; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _T_116; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_118; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [25:0] _T_120; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [25:0] _GEN_3; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_121; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_122; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_124; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [13:0] _GEN_4; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [14:0] _T_125; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire [7:0] _T_130; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  _T_139; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _T_142; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _T_143; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  _T_144; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire [5:0] _T_148; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _T_149; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _T_150; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _T_154; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _T_161; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _T_162; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _T_163; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _T_165; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  _T_170; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _T_172; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _T_174; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _T_175; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _T_177; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _T_178; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [8:0] _T_179; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] _T_181; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [8:0] _T_183; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [8:0] _T_185; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [8:0] _T_186; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [8:0] _T_188; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [8:0] _T_189; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [8:0] _T_191; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [8:0] _T_192; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [8:0] _T_193; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [8:0] _T_194; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [8:0] _T_195; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [8:0] _T_196; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [8:0] _T_197; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [8:0] _T_198; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_199; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _T_200; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [22:0] _T_201; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [22:0] _T_202; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [22:0] _T_204; // @[Bitwise.scala 72:12]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [9:0] _T_205; // @[Cat.scala 29:58]
  wire [1:0] _T_207; // @[Cat.scala 29:58]
  wire [2:0] _T_209; // @[Cat.scala 29:58]
  wire [29:0] RoundAnyRawFNToRecFN_3_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign sAdjustedExp = $signed(io_in_sExp) + $signed(-13'sh700); // @[RoundAnyRawFNToRecFN.scala 108:24]
  assign _T_5 = |io_in_sig[27:0]; // @[RoundAnyRawFNToRecFN.scala 115:60]
  assign adjustedSig = {io_in_sig[53:28],_T_5}; // @[Cat.scala 29:58]
  assign _T_8 = ~sAdjustedExp[8]; // @[primitives.scala 57:25]
  assign _T_10 = ~sAdjustedExp[7]; // @[primitives.scala 57:25]
  assign _T_12 = ~sAdjustedExp[6]; // @[primitives.scala 57:25]
  assign _T_13 = ~sAdjustedExp[5:0]; // @[primitives.scala 58:26]
  assign _T_14 = -65'sh10000000000000000 >>> _T_13; // @[primitives.scala 77:58]
  assign _T_20 = {{8'd0}, _T_14[57:50]}; // @[Bitwise.scala 103:31]
  assign _T_22 = {_T_14[49:42], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_24 = _T_22 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_25 = _T_20 | _T_24; // @[Bitwise.scala 103:39]
  assign _GEN_0 = {{4'd0}, _T_25[15:4]}; // @[Bitwise.scala 103:31]
  assign _T_30 = _GEN_0 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_32 = {_T_25[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_34 = _T_32 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_35 = _T_30 | _T_34; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{2'd0}, _T_35[15:2]}; // @[Bitwise.scala 103:31]
  assign _T_40 = _GEN_1 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_42 = {_T_35[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_44 = _T_42 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_45 = _T_40 | _T_44; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{1'd0}, _T_45[15:1]}; // @[Bitwise.scala 103:31]
  assign _T_50 = _GEN_2 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_52 = {_T_45[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_54 = _T_52 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_55 = _T_50 | _T_54; // @[Bitwise.scala 103:39]
  assign _T_72 = {_T_55,_T_14[58],_T_14[59],_T_14[60],_T_14[61],_T_14[62],_T_14[63]}; // @[Cat.scala 29:58]
  assign _T_74 = _T_12 ? 22'h0 : ~_T_72; // @[primitives.scala 74:21]
  assign _T_76 = {~_T_74,3'h7}; // @[Cat.scala 29:58]
  assign _T_86 = {_T_14[0],_T_14[1],_T_14[2]}; // @[Cat.scala 29:58]
  assign _T_87 = _T_12 ? _T_86 : 3'h0; // @[primitives.scala 61:24]
  assign _T_88 = _T_10 ? _T_76 : {{22'd0}, _T_87}; // @[primitives.scala 66:24]
  assign _T_89 = _T_8 ? _T_88 : 25'h0; // @[primitives.scala 61:24]
  assign _T_91 = {_T_89,2'h3}; // @[Cat.scala 29:58]
  assign _T_93 = {1'h0,_T_91[26:1]}; // @[Cat.scala 29:58]
  assign _T_95 = ~_T_93 & _T_91; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _T_96 = adjustedSig & _T_95; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_97 = |_T_96; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_98 = adjustedSig & _T_93; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_99 = |_T_98; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign _T_100 = _T_97 | _T_99; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_101 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_102 = _T_101 & _T_97; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_103 = roundMagUp & _T_100; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_104 = _T_102 | _T_103; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_105 = adjustedSig | _T_91; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_107 = _T_105[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_108 = roundingMode_near_even & _T_97; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_110 = _T_108 & ~_T_99; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_112 = _T_110 ? _T_91[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_114 = _T_107 & ~_T_112; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_116 = adjustedSig & ~_T_91; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_118 = roundingMode_odd & _T_100; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_120 = _T_118 ? _T_95[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_3 = {{1'd0}, _T_116[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_121 = _GEN_3 | _T_120; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_122 = _T_104 ? _T_114 : _T_121; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_124 = {1'b0,$signed(_T_122[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_4 = {{11{_T_124[2]}},_T_124}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_125 = $signed(sAdjustedExp) + $signed(_GEN_4); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_125[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = _T_122[22:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  assign _T_130 = _T_125[14:7]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_T_130) >= 8'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(_T_125) < 15'sh6b; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign _T_139 = |adjustedSig[1:0]; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign _T_142 = _T_101 & adjustedSig[1]; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _T_143 = roundMagUp & _T_139; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign _T_144 = _T_142 | _T_143; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign _T_148 = sAdjustedExp[13:8]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _T_149 = $signed(_T_148) <= 6'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _T_150 = _T_100 & _T_149; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _T_154 = _T_150 & _T_91[2]; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _T_161 = ~_T_91[3] & _T_122[24]; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _T_162 = _T_161 & _T_97; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _T_163 = _T_162 & _T_144; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _T_165 = _T_154 & ~_T_163; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _T_165; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | _T_100; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign _T_170 = ~isNaNOut & ~io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _T_170 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _T_172 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _T_172; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _T_101 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _T_174 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _T_175 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _T_174 & _T_175; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _T_177 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = io_in_isInf | _T_177; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _T_178 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _T_179 = _T_178 ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_181 = common_expOut & ~_T_179; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_183 = pegMinNonzeroMagOut ? 9'h194 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _T_185 = _T_181 & ~_T_183; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _T_186 = pegMaxFiniteMagOut ? 9'h80 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _T_188 = _T_185 & ~_T_186; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _T_189 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_191 = _T_188 & ~_T_189; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_192 = pegMinNonzeroMagOut ? 9'h6b : 9'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _T_193 = _T_191 | _T_192; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _T_194 = pegMaxFiniteMagOut ? 9'h17f : 9'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _T_195 = _T_193 | _T_194; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _T_196 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _T_197 = _T_195 | _T_196; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_198 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _T_197 | _T_198; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _T_199 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _T_200 = _T_199 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _T_201 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _T_202 = _T_200 ? _T_201 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_204 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0; // @[Bitwise.scala 72:12]
  assign fractOut = _T_202 | _T_204; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign _T_205 = {signOut,expOut}; // @[Cat.scala 29:58]
  assign _T_207 = {underflow,inexact}; // @[Cat.scala 29:58]
  assign _T_209 = {io_invalidExc,1'h0,overflow}; // @[Cat.scala 29:58]
  assign io_out = {_T_205,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_209,_T_207}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_3_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_3_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNToRaw_preMul_1(
  input  [1:0]   io_op,
  input  [64:0]  io_a,
  input  [64:0]  io_b,
  input  [64:0]  io_c,
  output [52:0]  io_mulAddA,
  output [52:0]  io_mulAddB,
  output [105:0] io_mulAddC,
  output         io_toPostMul_isSigNaNAny,
  output         io_toPostMul_isNaNAOrB,
  output         io_toPostMul_isInfA,
  output         io_toPostMul_isZeroA,
  output         io_toPostMul_isInfB,
  output         io_toPostMul_isZeroB,
  output         io_toPostMul_signProd,
  output         io_toPostMul_isNaNC,
  output         io_toPostMul_isInfC,
  output         io_toPostMul_isZeroC,
  output [12:0]  io_toPostMul_sExpSum,
  output         io_toPostMul_doSubMags,
  output         io_toPostMul_CIsDominant,
  output [5:0]   io_toPostMul_CDom_CAlignDist,
  output [54:0]  io_toPostMul_highAlignedSigC,
  output         io_toPostMul_bit0AlignedSigC,
  output [29:0]  io_covSum,
  output         metaAssert
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawA_sig; // @[Cat.scala 29:58]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawB_sig; // @[Cat.scala 29:58]
  wire  rawC_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_36; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawC_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawC_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawC_sig; // @[Cat.scala 29:58]
  wire  _T_48; // @[MulAddRecFN.scala 98:30]
  wire  signProd; // @[MulAddRecFN.scala 98:42]
  wire [13:0] _T_50; // @[MulAddRecFN.scala 101:19]
  wire [13:0] sExpAlignedProd; // @[MulAddRecFN.scala 101:32]
  wire  _T_53; // @[MulAddRecFN.scala 103:30]
  wire  doSubMags; // @[MulAddRecFN.scala 103:42]
  wire [13:0] _GEN_0; // @[MulAddRecFN.scala 107:42]
  wire [13:0] sNatCAlignDist; // @[MulAddRecFN.scala 107:42]
  wire [12:0] posNatCAlignDist; // @[MulAddRecFN.scala 108:42]
  wire  _T_57; // @[MulAddRecFN.scala 109:35]
  wire  _T_58; // @[MulAddRecFN.scala 109:69]
  wire  isMinCAlign; // @[MulAddRecFN.scala 109:50]
  wire  _T_60; // @[MulAddRecFN.scala 111:60]
  wire  _T_61; // @[MulAddRecFN.scala 111:39]
  wire  CIsDominant; // @[MulAddRecFN.scala 111:23]
  wire  _T_62; // @[MulAddRecFN.scala 115:34]
  wire [7:0] _T_64; // @[MulAddRecFN.scala 115:16]
  wire [7:0] CAlignDist; // @[MulAddRecFN.scala 113:12]
  wire [53:0] _T_66; // @[MulAddRecFN.scala 121:16]
  wire [110:0] _T_68; // @[Bitwise.scala 72:12]
  wire [164:0] _T_70; // @[MulAddRecFN.scala 123:11]
  wire [164:0] mainAlignedSigC; // @[MulAddRecFN.scala 123:17]
  wire  _T_74; // @[primitives.scala 121:54]
  wire  _T_76; // @[primitives.scala 121:54]
  wire  _T_78; // @[primitives.scala 121:54]
  wire  _T_80; // @[primitives.scala 121:54]
  wire  _T_82; // @[primitives.scala 121:54]
  wire  _T_84; // @[primitives.scala 121:54]
  wire  _T_86; // @[primitives.scala 121:54]
  wire  _T_88; // @[primitives.scala 121:54]
  wire  _T_90; // @[primitives.scala 121:54]
  wire  _T_92; // @[primitives.scala 121:54]
  wire  _T_94; // @[primitives.scala 121:54]
  wire  _T_96; // @[primitives.scala 121:54]
  wire  _T_98; // @[primitives.scala 121:54]
  wire  _T_100; // @[primitives.scala 124:57]
  wire [6:0] _T_106; // @[primitives.scala 125:20]
  wire [13:0] _T_113; // @[primitives.scala 125:20]
  wire [64:0] _T_115; // @[primitives.scala 77:58]
  wire [7:0] _T_121; // @[Bitwise.scala 103:31]
  wire [7:0] _T_123; // @[Bitwise.scala 103:65]
  wire [7:0] _T_125; // @[Bitwise.scala 103:75]
  wire [7:0] _T_126; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [7:0] _T_131; // @[Bitwise.scala 103:31]
  wire [7:0] _T_133; // @[Bitwise.scala 103:65]
  wire [7:0] _T_135; // @[Bitwise.scala 103:75]
  wire [7:0] _T_136; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [7:0] _T_141; // @[Bitwise.scala 103:31]
  wire [7:0] _T_143; // @[Bitwise.scala 103:65]
  wire [7:0] _T_145; // @[Bitwise.scala 103:75]
  wire [7:0] _T_146; // @[Bitwise.scala 103:39]
  wire [12:0] _T_160; // @[Cat.scala 29:58]
  wire [13:0] _GEN_3; // @[MulAddRecFN.scala 125:68]
  wire [13:0] _T_161; // @[MulAddRecFN.scala 125:68]
  wire  reduced4CExtra; // @[MulAddRecFN.scala 133:11]
  wire  _T_164; // @[MulAddRecFN.scala 137:39]
  wire  _T_166; // @[MulAddRecFN.scala 137:44]
  wire  _T_168; // @[MulAddRecFN.scala 138:39]
  wire  _T_169; // @[MulAddRecFN.scala 138:44]
  wire  _T_170; // @[MulAddRecFN.scala 136:16]
  wire [161:0] _T_171; // @[Cat.scala 29:58]
  wire [162:0] alignedSigC; // @[Cat.scala 29:58]
  wire  _T_175; // @[common.scala 81:46]
  wire  _T_178; // @[common.scala 81:46]
  wire  _T_179; // @[MulAddRecFN.scala 149:32]
  wire  _T_182; // @[common.scala 81:46]
  wire [13:0] _T_187; // @[MulAddRecFN.scala 161:53]
  wire [13:0] _T_188; // @[MulAddRecFN.scala 161:12]
  wire [29:0] MulAddRecFNToRaw_preMul_1_covSum;
  assign rawA_isZero = io_a[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_a[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_isNaN = _T_4 & io_a[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_sign = io_a[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_sExp = {1'b0,$signed(io_a[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_sig = {1'h0,~rawA_isZero,io_a[51:0]}; // @[Cat.scala 29:58]
  assign rawB_isZero = io_b[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_20 = io_b[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_isNaN = _T_20 & io_b[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_sign = io_b[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_sExp = {1'b0,$signed(io_b[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_sig = {1'h0,~rawB_isZero,io_b[51:0]}; // @[Cat.scala 29:58]
  assign rawC_isZero = io_c[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_36 = io_c[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawC_isNaN = _T_36 & io_c[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawC_sign = io_c[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawC_sExp = {1'b0,$signed(io_c[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawC_sig = {1'h0,~rawC_isZero,io_c[51:0]}; // @[Cat.scala 29:58]
  assign _T_48 = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30]
  assign signProd = _T_48 ^ io_op[1]; // @[MulAddRecFN.scala 98:42]
  assign _T_50 = $signed(rawA_sExp) + $signed(rawB_sExp); // @[MulAddRecFN.scala 101:19]
  assign sExpAlignedProd = $signed(_T_50) + -14'sh7c8; // @[MulAddRecFN.scala 101:32]
  assign _T_53 = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30]
  assign doSubMags = _T_53 ^ io_op[0]; // @[MulAddRecFN.scala 103:42]
  assign _GEN_0 = {{1{rawC_sExp[12]}},rawC_sExp}; // @[MulAddRecFN.scala 107:42]
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42]
  assign posNatCAlignDist = sNatCAlignDist[12:0]; // @[MulAddRecFN.scala 108:42]
  assign _T_57 = rawA_isZero | rawB_isZero; // @[MulAddRecFN.scala 109:35]
  assign _T_58 = $signed(sNatCAlignDist) < 14'sh0; // @[MulAddRecFN.scala 109:69]
  assign isMinCAlign = _T_57 | _T_58; // @[MulAddRecFN.scala 109:50]
  assign _T_60 = posNatCAlignDist <= 13'h35; // @[MulAddRecFN.scala 111:60]
  assign _T_61 = isMinCAlign | _T_60; // @[MulAddRecFN.scala 111:39]
  assign CIsDominant = ~rawC_isZero & _T_61; // @[MulAddRecFN.scala 111:23]
  assign _T_62 = posNatCAlignDist < 13'ha1; // @[MulAddRecFN.scala 115:34]
  assign _T_64 = _T_62 ? posNatCAlignDist[7:0] : 8'ha1; // @[MulAddRecFN.scala 115:16]
  assign CAlignDist = isMinCAlign ? 8'h0 : _T_64; // @[MulAddRecFN.scala 113:12]
  assign _T_66 = doSubMags ? ~rawC_sig : rawC_sig; // @[MulAddRecFN.scala 121:16]
  assign _T_68 = doSubMags ? 111'h7fffffffffffffffffffffffffff : 111'h0; // @[Bitwise.scala 72:12]
  assign _T_70 = {_T_66,_T_68}; // @[MulAddRecFN.scala 123:11]
  assign mainAlignedSigC = $signed(_T_70) >>> CAlignDist; // @[MulAddRecFN.scala 123:17]
  assign _T_74 = |rawC_sig[3:0]; // @[primitives.scala 121:54]
  assign _T_76 = |rawC_sig[7:4]; // @[primitives.scala 121:54]
  assign _T_78 = |rawC_sig[11:8]; // @[primitives.scala 121:54]
  assign _T_80 = |rawC_sig[15:12]; // @[primitives.scala 121:54]
  assign _T_82 = |rawC_sig[19:16]; // @[primitives.scala 121:54]
  assign _T_84 = |rawC_sig[23:20]; // @[primitives.scala 121:54]
  assign _T_86 = |rawC_sig[27:24]; // @[primitives.scala 121:54]
  assign _T_88 = |rawC_sig[31:28]; // @[primitives.scala 121:54]
  assign _T_90 = |rawC_sig[35:32]; // @[primitives.scala 121:54]
  assign _T_92 = |rawC_sig[39:36]; // @[primitives.scala 121:54]
  assign _T_94 = |rawC_sig[43:40]; // @[primitives.scala 121:54]
  assign _T_96 = |rawC_sig[47:44]; // @[primitives.scala 121:54]
  assign _T_98 = |rawC_sig[51:48]; // @[primitives.scala 121:54]
  assign _T_100 = |rawC_sig[53:52]; // @[primitives.scala 124:57]
  assign _T_106 = {_T_86,_T_84,_T_82,_T_80,_T_78,_T_76,_T_74}; // @[primitives.scala 125:20]
  assign _T_113 = {_T_100,_T_98,_T_96,_T_94,_T_92,_T_90,_T_88,_T_106}; // @[primitives.scala 125:20]
  assign _T_115 = -65'sh10000000000000000 >>> CAlignDist[7:2]; // @[primitives.scala 77:58]
  assign _T_121 = {{4'd0}, _T_115[31:28]}; // @[Bitwise.scala 103:31]
  assign _T_123 = {_T_115[27:24], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_125 = _T_123 & 8'hf0; // @[Bitwise.scala 103:75]
  assign _T_126 = _T_121 | _T_125; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{2'd0}, _T_126[7:2]}; // @[Bitwise.scala 103:31]
  assign _T_131 = _GEN_1 & 8'h33; // @[Bitwise.scala 103:31]
  assign _T_133 = {_T_126[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_135 = _T_133 & 8'hcc; // @[Bitwise.scala 103:75]
  assign _T_136 = _T_131 | _T_135; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{1'd0}, _T_136[7:1]}; // @[Bitwise.scala 103:31]
  assign _T_141 = _GEN_2 & 8'h55; // @[Bitwise.scala 103:31]
  assign _T_143 = {_T_136[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_145 = _T_143 & 8'haa; // @[Bitwise.scala 103:75]
  assign _T_146 = _T_141 | _T_145; // @[Bitwise.scala 103:39]
  assign _T_160 = {_T_146,_T_115[32],_T_115[33],_T_115[34],_T_115[35],_T_115[36]}; // @[Cat.scala 29:58]
  assign _GEN_3 = {{1'd0}, _T_160}; // @[MulAddRecFN.scala 125:68]
  assign _T_161 = _T_113 & _GEN_3; // @[MulAddRecFN.scala 125:68]
  assign reduced4CExtra = |_T_161; // @[MulAddRecFN.scala 133:11]
  assign _T_164 = &mainAlignedSigC[2:0]; // @[MulAddRecFN.scala 137:39]
  assign _T_166 = _T_164 & ~reduced4CExtra; // @[MulAddRecFN.scala 137:44]
  assign _T_168 = |mainAlignedSigC[2:0]; // @[MulAddRecFN.scala 138:39]
  assign _T_169 = _T_168 | reduced4CExtra; // @[MulAddRecFN.scala 138:44]
  assign _T_170 = doSubMags ? _T_166 : _T_169; // @[MulAddRecFN.scala 136:16]
  assign _T_171 = mainAlignedSigC[164:3]; // @[Cat.scala 29:58]
  assign alignedSigC = {_T_171,_T_170}; // @[Cat.scala 29:58]
  assign _T_175 = rawA_isNaN & ~rawA_sig[51]; // @[common.scala 81:46]
  assign _T_178 = rawB_isNaN & ~rawB_sig[51]; // @[common.scala 81:46]
  assign _T_179 = _T_175 | _T_178; // @[MulAddRecFN.scala 149:32]
  assign _T_182 = rawC_isNaN & ~rawC_sig[51]; // @[common.scala 81:46]
  assign _T_187 = $signed(sExpAlignedProd) - 14'sh35; // @[MulAddRecFN.scala 161:53]
  assign _T_188 = CIsDominant ? $signed({{1{rawC_sExp[12]}},rawC_sExp}) : $signed(_T_187); // @[MulAddRecFN.scala 161:12]
  assign io_mulAddA = rawA_sig[52:0]; // @[MulAddRecFN.scala 144:16]
  assign io_mulAddB = rawB_sig[52:0]; // @[MulAddRecFN.scala 145:16]
  assign io_mulAddC = alignedSigC[106:1]; // @[MulAddRecFN.scala 146:16]
  assign io_toPostMul_isSigNaNAny = _T_179 | _T_182; // @[MulAddRecFN.scala 148:30]
  assign io_toPostMul_isNaNAOrB = rawA_isNaN | rawB_isNaN; // @[MulAddRecFN.scala 151:28]
  assign io_toPostMul_isInfA = _T_4 & ~io_a[61]; // @[MulAddRecFN.scala 152:28]
  assign io_toPostMul_isZeroA = io_a[63:61] == 3'h0; // @[MulAddRecFN.scala 153:28]
  assign io_toPostMul_isInfB = _T_20 & ~io_b[61]; // @[MulAddRecFN.scala 154:28]
  assign io_toPostMul_isZeroB = io_b[63:61] == 3'h0; // @[MulAddRecFN.scala 155:28]
  assign io_toPostMul_signProd = _T_48 ^ io_op[1]; // @[MulAddRecFN.scala 156:28]
  assign io_toPostMul_isNaNC = _T_36 & io_c[61]; // @[MulAddRecFN.scala 157:28]
  assign io_toPostMul_isInfC = _T_36 & ~io_c[61]; // @[MulAddRecFN.scala 158:28]
  assign io_toPostMul_isZeroC = io_c[63:61] == 3'h0; // @[MulAddRecFN.scala 159:28]
  assign io_toPostMul_sExpSum = _T_188[12:0]; // @[MulAddRecFN.scala 160:28]
  assign io_toPostMul_doSubMags = _T_53 ^ io_op[0]; // @[MulAddRecFN.scala 162:28]
  assign io_toPostMul_CIsDominant = ~rawC_isZero & _T_61; // @[MulAddRecFN.scala 163:30]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[5:0]; // @[MulAddRecFN.scala 164:34]
  assign io_toPostMul_highAlignedSigC = alignedSigC[161:107]; // @[MulAddRecFN.scala 165:34]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:34]
  assign MulAddRecFNToRaw_preMul_1_covSum = 30'h0;
  assign io_covSum = MulAddRecFNToRaw_preMul_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNToRaw_postMul_1(
  input          io_fromPreMul_isSigNaNAny,
  input          io_fromPreMul_isNaNAOrB,
  input          io_fromPreMul_isInfA,
  input          io_fromPreMul_isZeroA,
  input          io_fromPreMul_isInfB,
  input          io_fromPreMul_isZeroB,
  input          io_fromPreMul_signProd,
  input          io_fromPreMul_isNaNC,
  input          io_fromPreMul_isInfC,
  input          io_fromPreMul_isZeroC,
  input  [12:0]  io_fromPreMul_sExpSum,
  input          io_fromPreMul_doSubMags,
  input          io_fromPreMul_CIsDominant,
  input  [5:0]   io_fromPreMul_CDom_CAlignDist,
  input  [54:0]  io_fromPreMul_highAlignedSigC,
  input          io_fromPreMul_bit0AlignedSigC,
  input  [106:0] io_mulAddResult,
  input  [2:0]   io_roundingMode,
  output         io_invalidExc,
  output         io_rawOut_isNaN,
  output         io_rawOut_isInf,
  output         io_rawOut_isZero,
  output         io_rawOut_sign,
  output [12:0]  io_rawOut_sExp,
  output [55:0]  io_rawOut_sig,
  output [29:0]  io_covSum,
  output         metaAssert
);
  wire  roundingMode_min; // @[MulAddRecFN.scala 188:45]
  wire  CDom_sign; // @[MulAddRecFN.scala 192:42]
  wire [54:0] _T_2; // @[MulAddRecFN.scala 195:47]
  wire [54:0] _T_3; // @[MulAddRecFN.scala 194:16]
  wire [161:0] sigSum; // @[Cat.scala 29:58]
  wire [1:0] _T_6; // @[MulAddRecFN.scala 205:69]
  wire [12:0] _GEN_0; // @[MulAddRecFN.scala 205:43]
  wire [12:0] CDom_sExp; // @[MulAddRecFN.scala 205:43]
  wire [107:0] _T_14; // @[Cat.scala 29:58]
  wire [107:0] CDom_absSigSum; // @[MulAddRecFN.scala 207:12]
  wire  _T_17; // @[MulAddRecFN.scala 217:36]
  wire  _T_19; // @[MulAddRecFN.scala 218:37]
  wire  CDom_absSigSumExtra; // @[MulAddRecFN.scala 216:12]
  wire [170:0] _GEN_1; // @[MulAddRecFN.scala 221:24]
  wire [170:0] _T_20; // @[MulAddRecFN.scala 221:24]
  wire [57:0] CDom_mainSig; // @[MulAddRecFN.scala 221:56]
  wire [54:0] _T_22; // @[MulAddRecFN.scala 224:53]
  wire  _T_25; // @[primitives.scala 121:54]
  wire  _T_27; // @[primitives.scala 121:54]
  wire  _T_29; // @[primitives.scala 121:54]
  wire  _T_31; // @[primitives.scala 121:54]
  wire  _T_33; // @[primitives.scala 121:54]
  wire  _T_35; // @[primitives.scala 121:54]
  wire  _T_37; // @[primitives.scala 121:54]
  wire  _T_39; // @[primitives.scala 121:54]
  wire  _T_41; // @[primitives.scala 121:54]
  wire  _T_43; // @[primitives.scala 121:54]
  wire  _T_45; // @[primitives.scala 121:54]
  wire  _T_47; // @[primitives.scala 121:54]
  wire  _T_49; // @[primitives.scala 121:54]
  wire  _T_51; // @[primitives.scala 124:57]
  wire [6:0] _T_57; // @[primitives.scala 125:20]
  wire [13:0] _T_64; // @[primitives.scala 125:20]
  wire [16:0] _T_67; // @[primitives.scala 77:58]
  wire [7:0] _T_73; // @[Bitwise.scala 103:31]
  wire [7:0] _T_75; // @[Bitwise.scala 103:65]
  wire [7:0] _T_77; // @[Bitwise.scala 103:75]
  wire [7:0] _T_78; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [7:0] _T_83; // @[Bitwise.scala 103:31]
  wire [7:0] _T_85; // @[Bitwise.scala 103:65]
  wire [7:0] _T_87; // @[Bitwise.scala 103:75]
  wire [7:0] _T_88; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_3; // @[Bitwise.scala 103:31]
  wire [7:0] _T_93; // @[Bitwise.scala 103:31]
  wire [7:0] _T_95; // @[Bitwise.scala 103:65]
  wire [7:0] _T_97; // @[Bitwise.scala 103:75]
  wire [7:0] _T_98; // @[Bitwise.scala 103:39]
  wire [12:0] _T_112; // @[Cat.scala 29:58]
  wire [13:0] _GEN_4; // @[MulAddRecFN.scala 224:72]
  wire [13:0] _T_113; // @[MulAddRecFN.scala 224:72]
  wire  CDom_reduced4SigExtra; // @[MulAddRecFN.scala 225:73]
  wire  _T_116; // @[MulAddRecFN.scala 228:32]
  wire  _T_117; // @[MulAddRecFN.scala 228:36]
  wire  _T_118; // @[MulAddRecFN.scala 228:61]
  wire [55:0] CDom_sig; // @[Cat.scala 29:58]
  wire  notCDom_signSigSum; // @[MulAddRecFN.scala 234:36]
  wire [108:0] _GEN_5; // @[MulAddRecFN.scala 238:41]
  wire [108:0] _T_123; // @[MulAddRecFN.scala 238:41]
  wire [108:0] notCDom_absSigSum; // @[MulAddRecFN.scala 236:12]
  wire  _T_126; // @[primitives.scala 104:54]
  wire  _T_128; // @[primitives.scala 104:54]
  wire  _T_130; // @[primitives.scala 104:54]
  wire  _T_132; // @[primitives.scala 104:54]
  wire  _T_134; // @[primitives.scala 104:54]
  wire  _T_136; // @[primitives.scala 104:54]
  wire  _T_138; // @[primitives.scala 104:54]
  wire  _T_140; // @[primitives.scala 104:54]
  wire  _T_142; // @[primitives.scala 104:54]
  wire  _T_144; // @[primitives.scala 104:54]
  wire  _T_146; // @[primitives.scala 104:54]
  wire  _T_148; // @[primitives.scala 104:54]
  wire  _T_150; // @[primitives.scala 104:54]
  wire  _T_152; // @[primitives.scala 104:54]
  wire  _T_154; // @[primitives.scala 104:54]
  wire  _T_156; // @[primitives.scala 104:54]
  wire  _T_158; // @[primitives.scala 104:54]
  wire  _T_160; // @[primitives.scala 104:54]
  wire  _T_162; // @[primitives.scala 104:54]
  wire  _T_164; // @[primitives.scala 104:54]
  wire  _T_166; // @[primitives.scala 104:54]
  wire  _T_168; // @[primitives.scala 104:54]
  wire  _T_170; // @[primitives.scala 104:54]
  wire  _T_172; // @[primitives.scala 104:54]
  wire  _T_174; // @[primitives.scala 104:54]
  wire  _T_176; // @[primitives.scala 104:54]
  wire  _T_178; // @[primitives.scala 104:54]
  wire  _T_180; // @[primitives.scala 104:54]
  wire  _T_182; // @[primitives.scala 104:54]
  wire  _T_184; // @[primitives.scala 104:54]
  wire  _T_186; // @[primitives.scala 104:54]
  wire  _T_188; // @[primitives.scala 104:54]
  wire  _T_190; // @[primitives.scala 104:54]
  wire  _T_192; // @[primitives.scala 104:54]
  wire  _T_194; // @[primitives.scala 104:54]
  wire  _T_196; // @[primitives.scala 104:54]
  wire  _T_198; // @[primitives.scala 104:54]
  wire  _T_200; // @[primitives.scala 104:54]
  wire  _T_202; // @[primitives.scala 104:54]
  wire  _T_204; // @[primitives.scala 104:54]
  wire  _T_206; // @[primitives.scala 104:54]
  wire  _T_208; // @[primitives.scala 104:54]
  wire  _T_210; // @[primitives.scala 104:54]
  wire  _T_212; // @[primitives.scala 104:54]
  wire  _T_214; // @[primitives.scala 104:54]
  wire  _T_216; // @[primitives.scala 104:54]
  wire  _T_218; // @[primitives.scala 104:54]
  wire  _T_220; // @[primitives.scala 104:54]
  wire  _T_222; // @[primitives.scala 104:54]
  wire  _T_224; // @[primitives.scala 104:54]
  wire  _T_226; // @[primitives.scala 104:54]
  wire  _T_228; // @[primitives.scala 104:54]
  wire  _T_230; // @[primitives.scala 104:54]
  wire  _T_232; // @[primitives.scala 104:54]
  wire  _T_234; // @[primitives.scala 107:57]
  wire [5:0] _T_239; // @[primitives.scala 108:20]
  wire [12:0] _T_246; // @[primitives.scala 108:20]
  wire [6:0] _T_252; // @[primitives.scala 108:20]
  wire [26:0] _T_260; // @[primitives.scala 108:20]
  wire [6:0] _T_266; // @[primitives.scala 108:20]
  wire [13:0] _T_273; // @[primitives.scala 108:20]
  wire [6:0] _T_279; // @[primitives.scala 108:20]
  wire [54:0] notCDom_reduced2AbsSigSum; // @[primitives.scala 108:20]
  wire [5:0] _T_343; // @[Mux.scala 47:69]
  wire [5:0] _T_344; // @[Mux.scala 47:69]
  wire [5:0] _T_345; // @[Mux.scala 47:69]
  wire [5:0] _T_346; // @[Mux.scala 47:69]
  wire [5:0] _T_347; // @[Mux.scala 47:69]
  wire [5:0] _T_348; // @[Mux.scala 47:69]
  wire [5:0] _T_349; // @[Mux.scala 47:69]
  wire [5:0] _T_350; // @[Mux.scala 47:69]
  wire [5:0] _T_351; // @[Mux.scala 47:69]
  wire [5:0] _T_352; // @[Mux.scala 47:69]
  wire [5:0] _T_353; // @[Mux.scala 47:69]
  wire [5:0] _T_354; // @[Mux.scala 47:69]
  wire [5:0] _T_355; // @[Mux.scala 47:69]
  wire [5:0] _T_356; // @[Mux.scala 47:69]
  wire [5:0] _T_357; // @[Mux.scala 47:69]
  wire [5:0] _T_358; // @[Mux.scala 47:69]
  wire [5:0] _T_359; // @[Mux.scala 47:69]
  wire [5:0] _T_360; // @[Mux.scala 47:69]
  wire [5:0] _T_361; // @[Mux.scala 47:69]
  wire [5:0] _T_362; // @[Mux.scala 47:69]
  wire [5:0] _T_363; // @[Mux.scala 47:69]
  wire [5:0] _T_364; // @[Mux.scala 47:69]
  wire [5:0] _T_365; // @[Mux.scala 47:69]
  wire [5:0] _T_366; // @[Mux.scala 47:69]
  wire [5:0] _T_367; // @[Mux.scala 47:69]
  wire [5:0] _T_368; // @[Mux.scala 47:69]
  wire [5:0] _T_369; // @[Mux.scala 47:69]
  wire [5:0] _T_370; // @[Mux.scala 47:69]
  wire [5:0] _T_371; // @[Mux.scala 47:69]
  wire [5:0] _T_372; // @[Mux.scala 47:69]
  wire [5:0] _T_373; // @[Mux.scala 47:69]
  wire [5:0] _T_374; // @[Mux.scala 47:69]
  wire [5:0] _T_375; // @[Mux.scala 47:69]
  wire [5:0] _T_376; // @[Mux.scala 47:69]
  wire [5:0] _T_377; // @[Mux.scala 47:69]
  wire [5:0] _T_378; // @[Mux.scala 47:69]
  wire [5:0] _T_379; // @[Mux.scala 47:69]
  wire [5:0] _T_380; // @[Mux.scala 47:69]
  wire [5:0] _T_381; // @[Mux.scala 47:69]
  wire [5:0] _T_382; // @[Mux.scala 47:69]
  wire [5:0] _T_383; // @[Mux.scala 47:69]
  wire [5:0] _T_384; // @[Mux.scala 47:69]
  wire [5:0] _T_385; // @[Mux.scala 47:69]
  wire [5:0] _T_386; // @[Mux.scala 47:69]
  wire [5:0] _T_387; // @[Mux.scala 47:69]
  wire [5:0] _T_388; // @[Mux.scala 47:69]
  wire [5:0] _T_389; // @[Mux.scala 47:69]
  wire [5:0] _T_390; // @[Mux.scala 47:69]
  wire [5:0] _T_391; // @[Mux.scala 47:69]
  wire [5:0] _T_392; // @[Mux.scala 47:69]
  wire [5:0] _T_393; // @[Mux.scala 47:69]
  wire [5:0] _T_394; // @[Mux.scala 47:69]
  wire [5:0] _T_395; // @[Mux.scala 47:69]
  wire [5:0] notCDom_normDistReduced2; // @[Mux.scala 47:69]
  wire [6:0] notCDom_nearNormDist; // @[MulAddRecFN.scala 242:56]
  wire [7:0] _T_396; // @[MulAddRecFN.scala 243:69]
  wire [12:0] _GEN_6; // @[MulAddRecFN.scala 243:46]
  wire [12:0] notCDom_sExp; // @[MulAddRecFN.scala 243:46]
  wire [235:0] _GEN_7; // @[MulAddRecFN.scala 245:27]
  wire [235:0] _T_399; // @[MulAddRecFN.scala 245:27]
  wire [57:0] notCDom_mainSig; // @[MulAddRecFN.scala 245:50]
  wire  _T_404; // @[primitives.scala 104:54]
  wire  _T_406; // @[primitives.scala 104:54]
  wire  _T_408; // @[primitives.scala 104:54]
  wire  _T_410; // @[primitives.scala 104:54]
  wire  _T_412; // @[primitives.scala 104:54]
  wire  _T_414; // @[primitives.scala 104:54]
  wire  _T_416; // @[primitives.scala 104:54]
  wire  _T_418; // @[primitives.scala 104:54]
  wire  _T_420; // @[primitives.scala 104:54]
  wire  _T_422; // @[primitives.scala 104:54]
  wire  _T_424; // @[primitives.scala 104:54]
  wire  _T_426; // @[primitives.scala 104:54]
  wire  _T_428; // @[primitives.scala 104:54]
  wire  _T_430; // @[primitives.scala 107:57]
  wire [6:0] _T_436; // @[primitives.scala 108:20]
  wire [13:0] _T_443; // @[primitives.scala 108:20]
  wire [32:0] _T_446; // @[primitives.scala 77:58]
  wire [7:0] _T_452; // @[Bitwise.scala 103:31]
  wire [7:0] _T_454; // @[Bitwise.scala 103:65]
  wire [7:0] _T_456; // @[Bitwise.scala 103:75]
  wire [7:0] _T_457; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_8; // @[Bitwise.scala 103:31]
  wire [7:0] _T_462; // @[Bitwise.scala 103:31]
  wire [7:0] _T_464; // @[Bitwise.scala 103:65]
  wire [7:0] _T_466; // @[Bitwise.scala 103:75]
  wire [7:0] _T_467; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_9; // @[Bitwise.scala 103:31]
  wire [7:0] _T_472; // @[Bitwise.scala 103:31]
  wire [7:0] _T_474; // @[Bitwise.scala 103:65]
  wire [7:0] _T_476; // @[Bitwise.scala 103:75]
  wire [7:0] _T_477; // @[Bitwise.scala 103:39]
  wire [12:0] _T_491; // @[Cat.scala 29:58]
  wire [13:0] _GEN_10; // @[MulAddRecFN.scala 249:78]
  wire [13:0] _T_492; // @[MulAddRecFN.scala 249:78]
  wire  notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 251:11]
  wire  _T_495; // @[MulAddRecFN.scala 254:35]
  wire  _T_496; // @[MulAddRecFN.scala 254:39]
  wire [55:0] notCDom_sig; // @[Cat.scala 29:58]
  wire  notCDom_completeCancellation; // @[MulAddRecFN.scala 257:50]
  wire  _T_498; // @[MulAddRecFN.scala 261:36]
  wire  notCDom_sign; // @[MulAddRecFN.scala 259:12]
  wire  notNaN_isInfProd; // @[MulAddRecFN.scala 266:49]
  wire  notNaN_isInfOut; // @[MulAddRecFN.scala 267:44]
  wire  _T_499; // @[MulAddRecFN.scala 269:32]
  wire  notNaN_addZeros; // @[MulAddRecFN.scala 269:58]
  wire  _T_500; // @[MulAddRecFN.scala 274:31]
  wire  _T_501; // @[MulAddRecFN.scala 273:35]
  wire  _T_502; // @[MulAddRecFN.scala 275:32]
  wire  _T_503; // @[MulAddRecFN.scala 274:57]
  wire  _T_506; // @[MulAddRecFN.scala 276:36]
  wire  _T_507; // @[MulAddRecFN.scala 277:61]
  wire  _T_508; // @[MulAddRecFN.scala 278:35]
  wire  _T_512; // @[MulAddRecFN.scala 285:42]
  wire  _T_514; // @[MulAddRecFN.scala 287:27]
  wire  _T_515; // @[MulAddRecFN.scala 288:31]
  wire  _T_516; // @[MulAddRecFN.scala 287:54]
  wire  _T_518; // @[MulAddRecFN.scala 289:26]
  wire  _T_519; // @[MulAddRecFN.scala 289:48]
  wire  _T_520; // @[MulAddRecFN.scala 290:36]
  wire  _T_521; // @[MulAddRecFN.scala 288:43]
  wire  _T_522; // @[MulAddRecFN.scala 291:26]
  wire  _T_523; // @[MulAddRecFN.scala 292:37]
  wire  _T_524; // @[MulAddRecFN.scala 291:46]
  wire  _T_525; // @[MulAddRecFN.scala 290:48]
  wire  _T_528; // @[MulAddRecFN.scala 293:28]
  wire  _T_529; // @[MulAddRecFN.scala 294:17]
  wire  _T_530; // @[MulAddRecFN.scala 293:49]
  wire [29:0] MulAddRecFNToRaw_postMul_1_covSum;
  assign roundingMode_min = io_roundingMode == 3'h2; // @[MulAddRecFN.scala 188:45]
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42]
  assign _T_2 = io_fromPreMul_highAlignedSigC + 55'h1; // @[MulAddRecFN.scala 195:47]
  assign _T_3 = io_mulAddResult[106] ? _T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16]
  assign sigSum = {_T_3,io_mulAddResult[105:0],io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 29:58]
  assign _T_6 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69]
  assign _GEN_0 = {{11{_T_6[1]}},_T_6}; // @[MulAddRecFN.scala 205:43]
  assign CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43]
  assign _T_14 = {1'h0,io_fromPreMul_highAlignedSigC[54:53],sigSum[159:55]}; // @[Cat.scala 29:58]
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? ~sigSum[161:54] : _T_14; // @[MulAddRecFN.scala 207:12]
  assign _T_17 = |~sigSum[53:1]; // @[MulAddRecFN.scala 217:36]
  assign _T_19 = |sigSum[54:1]; // @[MulAddRecFN.scala 218:37]
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_17 : _T_19; // @[MulAddRecFN.scala 216:12]
  assign _GEN_1 = {{63'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24]
  assign _T_20 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24]
  assign CDom_mainSig = _T_20[107:50]; // @[MulAddRecFN.scala 221:56]
  assign _T_22 = {CDom_absSigSum[52:0], 2'h0}; // @[MulAddRecFN.scala 224:53]
  assign _T_25 = |_T_22[3:0]; // @[primitives.scala 121:54]
  assign _T_27 = |_T_22[7:4]; // @[primitives.scala 121:54]
  assign _T_29 = |_T_22[11:8]; // @[primitives.scala 121:54]
  assign _T_31 = |_T_22[15:12]; // @[primitives.scala 121:54]
  assign _T_33 = |_T_22[19:16]; // @[primitives.scala 121:54]
  assign _T_35 = |_T_22[23:20]; // @[primitives.scala 121:54]
  assign _T_37 = |_T_22[27:24]; // @[primitives.scala 121:54]
  assign _T_39 = |_T_22[31:28]; // @[primitives.scala 121:54]
  assign _T_41 = |_T_22[35:32]; // @[primitives.scala 121:54]
  assign _T_43 = |_T_22[39:36]; // @[primitives.scala 121:54]
  assign _T_45 = |_T_22[43:40]; // @[primitives.scala 121:54]
  assign _T_47 = |_T_22[47:44]; // @[primitives.scala 121:54]
  assign _T_49 = |_T_22[51:48]; // @[primitives.scala 121:54]
  assign _T_51 = |_T_22[54:52]; // @[primitives.scala 124:57]
  assign _T_57 = {_T_37,_T_35,_T_33,_T_31,_T_29,_T_27,_T_25}; // @[primitives.scala 125:20]
  assign _T_64 = {_T_51,_T_49,_T_47,_T_45,_T_43,_T_41,_T_39,_T_57}; // @[primitives.scala 125:20]
  assign _T_67 = -17'sh10000 >>> ~io_fromPreMul_CDom_CAlignDist[5:2]; // @[primitives.scala 77:58]
  assign _T_73 = {{4'd0}, _T_67[8:5]}; // @[Bitwise.scala 103:31]
  assign _T_75 = {_T_67[4:1], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_77 = _T_75 & 8'hf0; // @[Bitwise.scala 103:75]
  assign _T_78 = _T_73 | _T_77; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{2'd0}, _T_78[7:2]}; // @[Bitwise.scala 103:31]
  assign _T_83 = _GEN_2 & 8'h33; // @[Bitwise.scala 103:31]
  assign _T_85 = {_T_78[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_87 = _T_85 & 8'hcc; // @[Bitwise.scala 103:75]
  assign _T_88 = _T_83 | _T_87; // @[Bitwise.scala 103:39]
  assign _GEN_3 = {{1'd0}, _T_88[7:1]}; // @[Bitwise.scala 103:31]
  assign _T_93 = _GEN_3 & 8'h55; // @[Bitwise.scala 103:31]
  assign _T_95 = {_T_88[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_97 = _T_95 & 8'haa; // @[Bitwise.scala 103:75]
  assign _T_98 = _T_93 | _T_97; // @[Bitwise.scala 103:39]
  assign _T_112 = {_T_98,_T_67[9],_T_67[10],_T_67[11],_T_67[12],_T_67[13]}; // @[Cat.scala 29:58]
  assign _GEN_4 = {{1'd0}, _T_112}; // @[MulAddRecFN.scala 224:72]
  assign _T_113 = _T_64 & _GEN_4; // @[MulAddRecFN.scala 224:72]
  assign CDom_reduced4SigExtra = |_T_113; // @[MulAddRecFN.scala 225:73]
  assign _T_116 = |CDom_mainSig[2:0]; // @[MulAddRecFN.scala 228:32]
  assign _T_117 = _T_116 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36]
  assign _T_118 = _T_117 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61]
  assign CDom_sig = {CDom_mainSig[57:3],_T_118}; // @[Cat.scala 29:58]
  assign notCDom_signSigSum = sigSum[109]; // @[MulAddRecFN.scala 234:36]
  assign _GEN_5 = {{108'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41]
  assign _T_123 = sigSum[108:0] + _GEN_5; // @[MulAddRecFN.scala 238:41]
  assign notCDom_absSigSum = notCDom_signSigSum ? ~sigSum[108:0] : _T_123; // @[MulAddRecFN.scala 236:12]
  assign _T_126 = |notCDom_absSigSum[1:0]; // @[primitives.scala 104:54]
  assign _T_128 = |notCDom_absSigSum[3:2]; // @[primitives.scala 104:54]
  assign _T_130 = |notCDom_absSigSum[5:4]; // @[primitives.scala 104:54]
  assign _T_132 = |notCDom_absSigSum[7:6]; // @[primitives.scala 104:54]
  assign _T_134 = |notCDom_absSigSum[9:8]; // @[primitives.scala 104:54]
  assign _T_136 = |notCDom_absSigSum[11:10]; // @[primitives.scala 104:54]
  assign _T_138 = |notCDom_absSigSum[13:12]; // @[primitives.scala 104:54]
  assign _T_140 = |notCDom_absSigSum[15:14]; // @[primitives.scala 104:54]
  assign _T_142 = |notCDom_absSigSum[17:16]; // @[primitives.scala 104:54]
  assign _T_144 = |notCDom_absSigSum[19:18]; // @[primitives.scala 104:54]
  assign _T_146 = |notCDom_absSigSum[21:20]; // @[primitives.scala 104:54]
  assign _T_148 = |notCDom_absSigSum[23:22]; // @[primitives.scala 104:54]
  assign _T_150 = |notCDom_absSigSum[25:24]; // @[primitives.scala 104:54]
  assign _T_152 = |notCDom_absSigSum[27:26]; // @[primitives.scala 104:54]
  assign _T_154 = |notCDom_absSigSum[29:28]; // @[primitives.scala 104:54]
  assign _T_156 = |notCDom_absSigSum[31:30]; // @[primitives.scala 104:54]
  assign _T_158 = |notCDom_absSigSum[33:32]; // @[primitives.scala 104:54]
  assign _T_160 = |notCDom_absSigSum[35:34]; // @[primitives.scala 104:54]
  assign _T_162 = |notCDom_absSigSum[37:36]; // @[primitives.scala 104:54]
  assign _T_164 = |notCDom_absSigSum[39:38]; // @[primitives.scala 104:54]
  assign _T_166 = |notCDom_absSigSum[41:40]; // @[primitives.scala 104:54]
  assign _T_168 = |notCDom_absSigSum[43:42]; // @[primitives.scala 104:54]
  assign _T_170 = |notCDom_absSigSum[45:44]; // @[primitives.scala 104:54]
  assign _T_172 = |notCDom_absSigSum[47:46]; // @[primitives.scala 104:54]
  assign _T_174 = |notCDom_absSigSum[49:48]; // @[primitives.scala 104:54]
  assign _T_176 = |notCDom_absSigSum[51:50]; // @[primitives.scala 104:54]
  assign _T_178 = |notCDom_absSigSum[53:52]; // @[primitives.scala 104:54]
  assign _T_180 = |notCDom_absSigSum[55:54]; // @[primitives.scala 104:54]
  assign _T_182 = |notCDom_absSigSum[57:56]; // @[primitives.scala 104:54]
  assign _T_184 = |notCDom_absSigSum[59:58]; // @[primitives.scala 104:54]
  assign _T_186 = |notCDom_absSigSum[61:60]; // @[primitives.scala 104:54]
  assign _T_188 = |notCDom_absSigSum[63:62]; // @[primitives.scala 104:54]
  assign _T_190 = |notCDom_absSigSum[65:64]; // @[primitives.scala 104:54]
  assign _T_192 = |notCDom_absSigSum[67:66]; // @[primitives.scala 104:54]
  assign _T_194 = |notCDom_absSigSum[69:68]; // @[primitives.scala 104:54]
  assign _T_196 = |notCDom_absSigSum[71:70]; // @[primitives.scala 104:54]
  assign _T_198 = |notCDom_absSigSum[73:72]; // @[primitives.scala 104:54]
  assign _T_200 = |notCDom_absSigSum[75:74]; // @[primitives.scala 104:54]
  assign _T_202 = |notCDom_absSigSum[77:76]; // @[primitives.scala 104:54]
  assign _T_204 = |notCDom_absSigSum[79:78]; // @[primitives.scala 104:54]
  assign _T_206 = |notCDom_absSigSum[81:80]; // @[primitives.scala 104:54]
  assign _T_208 = |notCDom_absSigSum[83:82]; // @[primitives.scala 104:54]
  assign _T_210 = |notCDom_absSigSum[85:84]; // @[primitives.scala 104:54]
  assign _T_212 = |notCDom_absSigSum[87:86]; // @[primitives.scala 104:54]
  assign _T_214 = |notCDom_absSigSum[89:88]; // @[primitives.scala 104:54]
  assign _T_216 = |notCDom_absSigSum[91:90]; // @[primitives.scala 104:54]
  assign _T_218 = |notCDom_absSigSum[93:92]; // @[primitives.scala 104:54]
  assign _T_220 = |notCDom_absSigSum[95:94]; // @[primitives.scala 104:54]
  assign _T_222 = |notCDom_absSigSum[97:96]; // @[primitives.scala 104:54]
  assign _T_224 = |notCDom_absSigSum[99:98]; // @[primitives.scala 104:54]
  assign _T_226 = |notCDom_absSigSum[101:100]; // @[primitives.scala 104:54]
  assign _T_228 = |notCDom_absSigSum[103:102]; // @[primitives.scala 104:54]
  assign _T_230 = |notCDom_absSigSum[105:104]; // @[primitives.scala 104:54]
  assign _T_232 = |notCDom_absSigSum[107:106]; // @[primitives.scala 104:54]
  assign _T_234 = |notCDom_absSigSum[108]; // @[primitives.scala 107:57]
  assign _T_239 = {_T_136,_T_134,_T_132,_T_130,_T_128,_T_126}; // @[primitives.scala 108:20]
  assign _T_246 = {_T_150,_T_148,_T_146,_T_144,_T_142,_T_140,_T_138,_T_239}; // @[primitives.scala 108:20]
  assign _T_252 = {_T_164,_T_162,_T_160,_T_158,_T_156,_T_154,_T_152}; // @[primitives.scala 108:20]
  assign _T_260 = {_T_178,_T_176,_T_174,_T_172,_T_170,_T_168,_T_166,_T_252,_T_246}; // @[primitives.scala 108:20]
  assign _T_266 = {_T_192,_T_190,_T_188,_T_186,_T_184,_T_182,_T_180}; // @[primitives.scala 108:20]
  assign _T_273 = {_T_206,_T_204,_T_202,_T_200,_T_198,_T_196,_T_194,_T_266}; // @[primitives.scala 108:20]
  assign _T_279 = {_T_220,_T_218,_T_216,_T_214,_T_212,_T_210,_T_208}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum = {_T_234,_T_232,_T_230,_T_228,_T_226,_T_224,_T_222,_T_279,_T_273,_T_260}; // @[primitives.scala 108:20]
  assign _T_343 = notCDom_reduced2AbsSigSum[1] ? 6'h35 : 6'h36; // @[Mux.scala 47:69]
  assign _T_344 = notCDom_reduced2AbsSigSum[2] ? 6'h34 : _T_343; // @[Mux.scala 47:69]
  assign _T_345 = notCDom_reduced2AbsSigSum[3] ? 6'h33 : _T_344; // @[Mux.scala 47:69]
  assign _T_346 = notCDom_reduced2AbsSigSum[4] ? 6'h32 : _T_345; // @[Mux.scala 47:69]
  assign _T_347 = notCDom_reduced2AbsSigSum[5] ? 6'h31 : _T_346; // @[Mux.scala 47:69]
  assign _T_348 = notCDom_reduced2AbsSigSum[6] ? 6'h30 : _T_347; // @[Mux.scala 47:69]
  assign _T_349 = notCDom_reduced2AbsSigSum[7] ? 6'h2f : _T_348; // @[Mux.scala 47:69]
  assign _T_350 = notCDom_reduced2AbsSigSum[8] ? 6'h2e : _T_349; // @[Mux.scala 47:69]
  assign _T_351 = notCDom_reduced2AbsSigSum[9] ? 6'h2d : _T_350; // @[Mux.scala 47:69]
  assign _T_352 = notCDom_reduced2AbsSigSum[10] ? 6'h2c : _T_351; // @[Mux.scala 47:69]
  assign _T_353 = notCDom_reduced2AbsSigSum[11] ? 6'h2b : _T_352; // @[Mux.scala 47:69]
  assign _T_354 = notCDom_reduced2AbsSigSum[12] ? 6'h2a : _T_353; // @[Mux.scala 47:69]
  assign _T_355 = notCDom_reduced2AbsSigSum[13] ? 6'h29 : _T_354; // @[Mux.scala 47:69]
  assign _T_356 = notCDom_reduced2AbsSigSum[14] ? 6'h28 : _T_355; // @[Mux.scala 47:69]
  assign _T_357 = notCDom_reduced2AbsSigSum[15] ? 6'h27 : _T_356; // @[Mux.scala 47:69]
  assign _T_358 = notCDom_reduced2AbsSigSum[16] ? 6'h26 : _T_357; // @[Mux.scala 47:69]
  assign _T_359 = notCDom_reduced2AbsSigSum[17] ? 6'h25 : _T_358; // @[Mux.scala 47:69]
  assign _T_360 = notCDom_reduced2AbsSigSum[18] ? 6'h24 : _T_359; // @[Mux.scala 47:69]
  assign _T_361 = notCDom_reduced2AbsSigSum[19] ? 6'h23 : _T_360; // @[Mux.scala 47:69]
  assign _T_362 = notCDom_reduced2AbsSigSum[20] ? 6'h22 : _T_361; // @[Mux.scala 47:69]
  assign _T_363 = notCDom_reduced2AbsSigSum[21] ? 6'h21 : _T_362; // @[Mux.scala 47:69]
  assign _T_364 = notCDom_reduced2AbsSigSum[22] ? 6'h20 : _T_363; // @[Mux.scala 47:69]
  assign _T_365 = notCDom_reduced2AbsSigSum[23] ? 6'h1f : _T_364; // @[Mux.scala 47:69]
  assign _T_366 = notCDom_reduced2AbsSigSum[24] ? 6'h1e : _T_365; // @[Mux.scala 47:69]
  assign _T_367 = notCDom_reduced2AbsSigSum[25] ? 6'h1d : _T_366; // @[Mux.scala 47:69]
  assign _T_368 = notCDom_reduced2AbsSigSum[26] ? 6'h1c : _T_367; // @[Mux.scala 47:69]
  assign _T_369 = notCDom_reduced2AbsSigSum[27] ? 6'h1b : _T_368; // @[Mux.scala 47:69]
  assign _T_370 = notCDom_reduced2AbsSigSum[28] ? 6'h1a : _T_369; // @[Mux.scala 47:69]
  assign _T_371 = notCDom_reduced2AbsSigSum[29] ? 6'h19 : _T_370; // @[Mux.scala 47:69]
  assign _T_372 = notCDom_reduced2AbsSigSum[30] ? 6'h18 : _T_371; // @[Mux.scala 47:69]
  assign _T_373 = notCDom_reduced2AbsSigSum[31] ? 6'h17 : _T_372; // @[Mux.scala 47:69]
  assign _T_374 = notCDom_reduced2AbsSigSum[32] ? 6'h16 : _T_373; // @[Mux.scala 47:69]
  assign _T_375 = notCDom_reduced2AbsSigSum[33] ? 6'h15 : _T_374; // @[Mux.scala 47:69]
  assign _T_376 = notCDom_reduced2AbsSigSum[34] ? 6'h14 : _T_375; // @[Mux.scala 47:69]
  assign _T_377 = notCDom_reduced2AbsSigSum[35] ? 6'h13 : _T_376; // @[Mux.scala 47:69]
  assign _T_378 = notCDom_reduced2AbsSigSum[36] ? 6'h12 : _T_377; // @[Mux.scala 47:69]
  assign _T_379 = notCDom_reduced2AbsSigSum[37] ? 6'h11 : _T_378; // @[Mux.scala 47:69]
  assign _T_380 = notCDom_reduced2AbsSigSum[38] ? 6'h10 : _T_379; // @[Mux.scala 47:69]
  assign _T_381 = notCDom_reduced2AbsSigSum[39] ? 6'hf : _T_380; // @[Mux.scala 47:69]
  assign _T_382 = notCDom_reduced2AbsSigSum[40] ? 6'he : _T_381; // @[Mux.scala 47:69]
  assign _T_383 = notCDom_reduced2AbsSigSum[41] ? 6'hd : _T_382; // @[Mux.scala 47:69]
  assign _T_384 = notCDom_reduced2AbsSigSum[42] ? 6'hc : _T_383; // @[Mux.scala 47:69]
  assign _T_385 = notCDom_reduced2AbsSigSum[43] ? 6'hb : _T_384; // @[Mux.scala 47:69]
  assign _T_386 = notCDom_reduced2AbsSigSum[44] ? 6'ha : _T_385; // @[Mux.scala 47:69]
  assign _T_387 = notCDom_reduced2AbsSigSum[45] ? 6'h9 : _T_386; // @[Mux.scala 47:69]
  assign _T_388 = notCDom_reduced2AbsSigSum[46] ? 6'h8 : _T_387; // @[Mux.scala 47:69]
  assign _T_389 = notCDom_reduced2AbsSigSum[47] ? 6'h7 : _T_388; // @[Mux.scala 47:69]
  assign _T_390 = notCDom_reduced2AbsSigSum[48] ? 6'h6 : _T_389; // @[Mux.scala 47:69]
  assign _T_391 = notCDom_reduced2AbsSigSum[49] ? 6'h5 : _T_390; // @[Mux.scala 47:69]
  assign _T_392 = notCDom_reduced2AbsSigSum[50] ? 6'h4 : _T_391; // @[Mux.scala 47:69]
  assign _T_393 = notCDom_reduced2AbsSigSum[51] ? 6'h3 : _T_392; // @[Mux.scala 47:69]
  assign _T_394 = notCDom_reduced2AbsSigSum[52] ? 6'h2 : _T_393; // @[Mux.scala 47:69]
  assign _T_395 = notCDom_reduced2AbsSigSum[53] ? 6'h1 : _T_394; // @[Mux.scala 47:69]
  assign notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[54] ? 6'h0 : _T_395; // @[Mux.scala 47:69]
  assign notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56]
  assign _T_396 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69]
  assign _GEN_6 = {{5{_T_396[7]}},_T_396}; // @[MulAddRecFN.scala 243:46]
  assign notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_6); // @[MulAddRecFN.scala 243:46]
  assign _GEN_7 = {{127'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27]
  assign _T_399 = _GEN_7 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27]
  assign notCDom_mainSig = _T_399[109:52]; // @[MulAddRecFN.scala 245:50]
  assign _T_404 = |notCDom_reduced2AbsSigSum[1:0]; // @[primitives.scala 104:54]
  assign _T_406 = |notCDom_reduced2AbsSigSum[3:2]; // @[primitives.scala 104:54]
  assign _T_408 = |notCDom_reduced2AbsSigSum[5:4]; // @[primitives.scala 104:54]
  assign _T_410 = |notCDom_reduced2AbsSigSum[7:6]; // @[primitives.scala 104:54]
  assign _T_412 = |notCDom_reduced2AbsSigSum[9:8]; // @[primitives.scala 104:54]
  assign _T_414 = |notCDom_reduced2AbsSigSum[11:10]; // @[primitives.scala 104:54]
  assign _T_416 = |notCDom_reduced2AbsSigSum[13:12]; // @[primitives.scala 104:54]
  assign _T_418 = |notCDom_reduced2AbsSigSum[15:14]; // @[primitives.scala 104:54]
  assign _T_420 = |notCDom_reduced2AbsSigSum[17:16]; // @[primitives.scala 104:54]
  assign _T_422 = |notCDom_reduced2AbsSigSum[19:18]; // @[primitives.scala 104:54]
  assign _T_424 = |notCDom_reduced2AbsSigSum[21:20]; // @[primitives.scala 104:54]
  assign _T_426 = |notCDom_reduced2AbsSigSum[23:22]; // @[primitives.scala 104:54]
  assign _T_428 = |notCDom_reduced2AbsSigSum[25:24]; // @[primitives.scala 104:54]
  assign _T_430 = |notCDom_reduced2AbsSigSum[26]; // @[primitives.scala 107:57]
  assign _T_436 = {_T_416,_T_414,_T_412,_T_410,_T_408,_T_406,_T_404}; // @[primitives.scala 108:20]
  assign _T_443 = {_T_430,_T_428,_T_426,_T_424,_T_422,_T_420,_T_418,_T_436}; // @[primitives.scala 108:20]
  assign _T_446 = -33'sh100000000 >>> ~notCDom_normDistReduced2[5:1]; // @[primitives.scala 77:58]
  assign _T_452 = {{4'd0}, _T_446[8:5]}; // @[Bitwise.scala 103:31]
  assign _T_454 = {_T_446[4:1], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_456 = _T_454 & 8'hf0; // @[Bitwise.scala 103:75]
  assign _T_457 = _T_452 | _T_456; // @[Bitwise.scala 103:39]
  assign _GEN_8 = {{2'd0}, _T_457[7:2]}; // @[Bitwise.scala 103:31]
  assign _T_462 = _GEN_8 & 8'h33; // @[Bitwise.scala 103:31]
  assign _T_464 = {_T_457[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_466 = _T_464 & 8'hcc; // @[Bitwise.scala 103:75]
  assign _T_467 = _T_462 | _T_466; // @[Bitwise.scala 103:39]
  assign _GEN_9 = {{1'd0}, _T_467[7:1]}; // @[Bitwise.scala 103:31]
  assign _T_472 = _GEN_9 & 8'h55; // @[Bitwise.scala 103:31]
  assign _T_474 = {_T_467[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_476 = _T_474 & 8'haa; // @[Bitwise.scala 103:75]
  assign _T_477 = _T_472 | _T_476; // @[Bitwise.scala 103:39]
  assign _T_491 = {_T_477,_T_446[9],_T_446[10],_T_446[11],_T_446[12],_T_446[13]}; // @[Cat.scala 29:58]
  assign _GEN_10 = {{1'd0}, _T_491}; // @[MulAddRecFN.scala 249:78]
  assign _T_492 = _T_443 & _GEN_10; // @[MulAddRecFN.scala 249:78]
  assign notCDom_reduced4SigExtra = |_T_492; // @[MulAddRecFN.scala 251:11]
  assign _T_495 = |notCDom_mainSig[2:0]; // @[MulAddRecFN.scala 254:35]
  assign _T_496 = _T_495 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39]
  assign notCDom_sig = {notCDom_mainSig[57:3],_T_496}; // @[Cat.scala 29:58]
  assign notCDom_completeCancellation = notCDom_sig[55:54] == 2'h0; // @[MulAddRecFN.scala 257:50]
  assign _T_498 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36]
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _T_498; // @[MulAddRecFN.scala 259:12]
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49]
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  assign _T_499 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32]
  assign notNaN_addZeros = _T_499 & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58]
  assign _T_500 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31]
  assign _T_501 = io_fromPreMul_isSigNaNAny | _T_500; // @[MulAddRecFN.scala 273:35]
  assign _T_502 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32]
  assign _T_503 = _T_501 | _T_502; // @[MulAddRecFN.scala 274:57]
  assign _T_506 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36]
  assign _T_507 = _T_506 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61]
  assign _T_508 = _T_507 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35]
  assign _T_512 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42]
  assign _T_514 = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27]
  assign _T_515 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31]
  assign _T_516 = _T_514 | _T_515; // @[MulAddRecFN.scala 287:54]
  assign _T_518 = notNaN_addZeros & ~roundingMode_min; // @[MulAddRecFN.scala 289:26]
  assign _T_519 = _T_518 & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48]
  assign _T_520 = _T_519 & CDom_sign; // @[MulAddRecFN.scala 290:36]
  assign _T_521 = _T_516 | _T_520; // @[MulAddRecFN.scala 288:43]
  assign _T_522 = notNaN_addZeros & roundingMode_min; // @[MulAddRecFN.scala 291:26]
  assign _T_523 = io_fromPreMul_signProd | CDom_sign; // @[MulAddRecFN.scala 292:37]
  assign _T_524 = _T_522 & _T_523; // @[MulAddRecFN.scala 291:46]
  assign _T_525 = _T_521 | _T_524; // @[MulAddRecFN.scala 290:48]
  assign _T_528 = ~notNaN_isInfOut & ~notNaN_addZeros; // @[MulAddRecFN.scala 293:28]
  assign _T_529 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17]
  assign _T_530 = _T_528 & _T_529; // @[MulAddRecFN.scala 293:49]
  assign io_invalidExc = _T_503 | _T_508; // @[MulAddRecFN.scala 272:19]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21]
  assign io_rawOut_isZero = notNaN_addZeros | _T_512; // @[MulAddRecFN.scala 283:22]
  assign io_rawOut_sign = _T_525 | _T_530; // @[MulAddRecFN.scala 286:20]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19]
  assign MulAddRecFNToRaw_postMul_1_covSum = 30'h0;
  assign io_covSum = MulAddRecFNToRaw_postMul_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module DivSqrtRawFN_small(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [9:0]  io_a_sExp,
  input  [24:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [9:0]  io_b_sExp,
  input  [24:0] io_b_sig,
  input  [2:0]  io_roundingMode,
  output        io_rawOutValid_div,
  output        io_rawOutValid_sqrt,
  output [2:0]  io_roundingModeOut,
  output        io_invalidExc,
  output        io_infiniteExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [26:0] cycleNum; // @[DivSqrtRecFN_small.scala 223:33]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[DivSqrtRecFN_small.scala 225:29]
  reg [31:0] _RAND_1;
  reg  majorExc_Z; // @[DivSqrtRecFN_small.scala 226:29]
  reg [31:0] _RAND_2;
  reg  isNaN_Z; // @[DivSqrtRecFN_small.scala 228:29]
  reg [31:0] _RAND_3;
  reg  isInf_Z; // @[DivSqrtRecFN_small.scala 229:29]
  reg [31:0] _RAND_4;
  reg  isZero_Z; // @[DivSqrtRecFN_small.scala 230:29]
  reg [31:0] _RAND_5;
  reg  sign_Z; // @[DivSqrtRecFN_small.scala 231:29]
  reg [31:0] _RAND_6;
  reg [9:0] sExp_Z; // @[DivSqrtRecFN_small.scala 232:29]
  reg [31:0] _RAND_7;
  reg [22:0] fractB_Z; // @[DivSqrtRecFN_small.scala 233:29]
  reg [31:0] _RAND_8;
  reg [2:0] roundingMode_Z; // @[DivSqrtRecFN_small.scala 234:29]
  reg [31:0] _RAND_9;
  reg [25:0] rem_Z; // @[DivSqrtRecFN_small.scala 240:29]
  reg [31:0] _RAND_10;
  reg  notZeroRem_Z; // @[DivSqrtRecFN_small.scala 241:29]
  reg [31:0] _RAND_11;
  reg [25:0] sigX_Z; // @[DivSqrtRecFN_small.scala 242:29]
  reg [31:0] _RAND_12;
  wire  _T; // @[DivSqrtRecFN_small.scala 251:24]
  wire  _T_1; // @[DivSqrtRecFN_small.scala 251:59]
  wire  notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 251:42]
  wire  _T_4; // @[DivSqrtRecFN_small.scala 253:24]
  wire  notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 253:43]
  wire  _T_7; // @[common.scala 81:46]
  wire  _T_8; // @[DivSqrtRecFN_small.scala 256:38]
  wire  _T_14; // @[common.scala 81:46]
  wire  _T_15; // @[DivSqrtRecFN_small.scala 257:38]
  wire  _T_16; // @[DivSqrtRecFN_small.scala 257:66]
  wire  _T_19; // @[DivSqrtRecFN_small.scala 259:33]
  wire  _T_20; // @[DivSqrtRecFN_small.scala 259:51]
  wire  _T_21; // @[DivSqrtRecFN_small.scala 258:46]
  wire  _T_22; // @[DivSqrtRecFN_small.scala 263:26]
  wire  _T_23; // @[DivSqrtRecFN_small.scala 264:26]
  wire  _T_24; // @[DivSqrtRecFN_small.scala 264:42]
  wire  _T_25; // @[DivSqrtRecFN_small.scala 266:63]
  wire  _T_26; // @[DivSqrtRecFN_small.scala 267:64]
  wire  _T_28; // @[DivSqrtRecFN_small.scala 268:45]
  wire  sign_S; // @[DivSqrtRecFN_small.scala 268:30]
  wire  _T_29; // @[DivSqrtRecFN_small.scala 270:39]
  wire  specialCaseA_S; // @[DivSqrtRecFN_small.scala 270:55]
  wire  _T_30; // @[DivSqrtRecFN_small.scala 271:39]
  wire  specialCaseB_S; // @[DivSqrtRecFN_small.scala 271:55]
  wire  normalCase_S_div; // @[DivSqrtRecFN_small.scala 272:45]
  wire  normalCase_S_sqrt; // @[DivSqrtRecFN_small.scala 273:46]
  wire  normalCase_S; // @[DivSqrtRecFN_small.scala 274:27]
  wire [8:0] _T_39; // @[DivSqrtRecFN_small.scala 278:71]
  wire [9:0] _GEN_13; // @[DivSqrtRecFN_small.scala 277:21]
  wire [10:0] sExpQuot_S_div; // @[DivSqrtRecFN_small.scala 277:21]
  wire  _T_40; // @[DivSqrtRecFN_small.scala 281:48]
  wire [3:0] _T_42; // @[DivSqrtRecFN_small.scala 281:16]
  wire [9:0] sSatExpQuot_S_div; // @[DivSqrtRecFN_small.scala 286:11]
  wire  evenSqrt_S; // @[DivSqrtRecFN_small.scala 288:32]
  wire  oddSqrt_S; // @[DivSqrtRecFN_small.scala 289:32]
  wire  idle; // @[DivSqrtRecFN_small.scala 293:24]
  wire  inReady; // @[DivSqrtRecFN_small.scala 294:24]
  wire  entering; // @[DivSqrtRecFN_small.scala 295:28]
  wire  entering_normalCase; // @[DivSqrtRecFN_small.scala 296:40]
  wire  skipCycle2; // @[DivSqrtRecFN_small.scala 298:34]
  wire  _T_52; // @[DivSqrtRecFN_small.scala 300:18]
  wire  _T_54; // @[DivSqrtRecFN_small.scala 302:26]
  wire [1:0] _T_55; // @[DivSqrtRecFN_small.scala 302:16]
  wire [25:0] _T_57; // @[DivSqrtRecFN_small.scala 305:24]
  wire [26:0] _T_58; // @[DivSqrtRecFN_small.scala 304:20]
  wire [26:0] _T_59; // @[DivSqrtRecFN_small.scala 303:16]
  wire [26:0] _GEN_14; // @[DivSqrtRecFN_small.scala 302:59]
  wire [26:0] _T_60; // @[DivSqrtRecFN_small.scala 302:59]
  wire  _T_63; // @[DivSqrtRecFN_small.scala 310:28]
  wire [25:0] _T_65; // @[DivSqrtRecFN_small.scala 310:16]
  wire [26:0] _GEN_15; // @[DivSqrtRecFN_small.scala 309:15]
  wire [26:0] _T_66; // @[DivSqrtRecFN_small.scala 309:15]
  wire [1:0] _T_67; // @[DivSqrtRecFN_small.scala 311:16]
  wire [26:0] _GEN_16; // @[DivSqrtRecFN_small.scala 310:63]
  wire [26:0] _T_68; // @[DivSqrtRecFN_small.scala 310:63]
  wire [8:0] _T_69; // @[DivSqrtRecFN_small.scala 329:29]
  wire [9:0] _T_70; // @[DivSqrtRecFN_small.scala 329:34]
  wire  _T_73; // @[DivSqrtRecFN_small.scala 334:31]
  wire  _T_76; // @[DivSqrtRecFN_small.scala 341:21]
  wire [25:0] _T_77; // @[DivSqrtRecFN_small.scala 341:47]
  wire [25:0] _T_78; // @[DivSqrtRecFN_small.scala 341:12]
  wire  _T_79; // @[DivSqrtRecFN_small.scala 342:21]
  wire [1:0] _T_82; // @[DivSqrtRecFN_small.scala 343:56]
  wire [24:0] _T_84; // @[DivSqrtRecFN_small.scala 344:44]
  wire [26:0] _T_85; // @[Cat.scala 29:58]
  wire [26:0] _T_86; // @[DivSqrtRecFN_small.scala 342:12]
  wire [26:0] _GEN_17; // @[DivSqrtRecFN_small.scala 341:57]
  wire [26:0] _T_87; // @[DivSqrtRecFN_small.scala 341:57]
  wire [26:0] _T_89; // @[DivSqrtRecFN_small.scala 348:29]
  wire [26:0] _T_90; // @[DivSqrtRecFN_small.scala 348:12]
  wire [26:0] rem; // @[DivSqrtRecFN_small.scala 347:11]
  wire [24:0] bitMask; // @[DivSqrtRecFN_small.scala 349:27]
  wire  _T_92; // @[DivSqrtRecFN_small.scala 351:21]
  wire [25:0] _T_93; // @[DivSqrtRecFN_small.scala 351:47]
  wire [25:0] _T_94; // @[DivSqrtRecFN_small.scala 351:12]
  wire  _T_95; // @[DivSqrtRecFN_small.scala 352:21]
  wire [24:0] _T_96; // @[DivSqrtRecFN_small.scala 352:12]
  wire [25:0] _GEN_18; // @[DivSqrtRecFN_small.scala 351:73]
  wire [25:0] _T_97; // @[DivSqrtRecFN_small.scala 351:73]
  wire [25:0] _T_99; // @[DivSqrtRecFN_small.scala 353:12]
  wire [25:0] _T_100; // @[DivSqrtRecFN_small.scala 352:73]
  wire  _T_103; // @[DivSqrtRecFN_small.scala 354:23]
  wire [23:0] _T_104; // @[Cat.scala 29:58]
  wire [24:0] _T_105; // @[DivSqrtRecFN_small.scala 354:56]
  wire [24:0] _T_106; // @[DivSqrtRecFN_small.scala 354:12]
  wire [25:0] _GEN_19; // @[DivSqrtRecFN_small.scala 353:73]
  wire [25:0] _T_107; // @[DivSqrtRecFN_small.scala 353:73]
  wire  _T_109; // @[DivSqrtRecFN_small.scala 355:23]
  wire [26:0] _T_110; // @[DivSqrtRecFN_small.scala 355:44]
  wire [26:0] _GEN_20; // @[DivSqrtRecFN_small.scala 355:48]
  wire [26:0] _T_111; // @[DivSqrtRecFN_small.scala 355:48]
  wire [26:0] _T_112; // @[DivSqrtRecFN_small.scala 355:12]
  wire [26:0] _GEN_21; // @[DivSqrtRecFN_small.scala 354:73]
  wire [26:0] trialTerm; // @[DivSqrtRecFN_small.scala 354:73]
  wire [27:0] _T_113; // @[DivSqrtRecFN_small.scala 356:24]
  wire [27:0] _T_114; // @[DivSqrtRecFN_small.scala 356:41]
  wire [27:0] trialRem; // @[DivSqrtRecFN_small.scala 356:29]
  wire  newBit; // @[DivSqrtRecFN_small.scala 357:23]
  wire  _T_118; // @[DivSqrtRecFN_small.scala 359:41]
  wire  _T_120; // @[DivSqrtRecFN_small.scala 359:31]
  wire [27:0] _T_121; // @[DivSqrtRecFN_small.scala 360:39]
  wire [27:0] _T_122; // @[DivSqrtRecFN_small.scala 360:21]
  wire [27:0] _GEN_10; // @[DivSqrtRecFN_small.scala 359:58]
  wire  _T_124; // @[DivSqrtRecFN_small.scala 362:45]
  wire  _T_125; // @[DivSqrtRecFN_small.scala 362:31]
  wire  _T_126; // @[DivSqrtRecFN_small.scala 363:35]
  wire [25:0] _T_129; // @[DivSqrtRecFN_small.scala 365:47]
  wire [25:0] _T_130; // @[DivSqrtRecFN_small.scala 365:16]
  wire  _T_131; // @[DivSqrtRecFN_small.scala 366:25]
  wire [24:0] _T_132; // @[DivSqrtRecFN_small.scala 366:16]
  wire [25:0] _GEN_22; // @[DivSqrtRecFN_small.scala 365:71]
  wire [25:0] _T_133; // @[DivSqrtRecFN_small.scala 365:71]
  wire [23:0] _T_135; // @[DivSqrtRecFN_small.scala 367:47]
  wire [23:0] _T_136; // @[DivSqrtRecFN_small.scala 367:16]
  wire [25:0] _GEN_23; // @[DivSqrtRecFN_small.scala 366:71]
  wire [25:0] _T_137; // @[DivSqrtRecFN_small.scala 366:71]
  wire [25:0] _GEN_24; // @[DivSqrtRecFN_small.scala 368:48]
  wire [25:0] _T_139; // @[DivSqrtRecFN_small.scala 368:48]
  wire [25:0] _T_140; // @[DivSqrtRecFN_small.scala 368:16]
  wire [25:0] _T_141; // @[DivSqrtRecFN_small.scala 367:71]
  wire [26:0] _GEN_25; // @[DivSqrtRecFN_small.scala 385:35]
  reg [4:0] DivSqrtRawFN_small_state; // @[Register tracking DivSqrtRawFN_small state]
  reg [31:0] _RAND_13;
  reg  DivSqrtRawFN_small_cov [0:31]; // @[Coverage map for DivSqrtRawFN_small]
  reg [31:0] _RAND_14;
  wire  DivSqrtRawFN_small_cov_read_data; // @[Coverage map for DivSqrtRawFN_small]
  wire [4:0] DivSqrtRawFN_small_cov_read_addr; // @[Coverage map for DivSqrtRawFN_small]
  wire  DivSqrtRawFN_small_cov_write_data; // @[Coverage map for DivSqrtRawFN_small]
  wire [4:0] DivSqrtRawFN_small_cov_write_addr; // @[Coverage map for DivSqrtRawFN_small]
  wire  DivSqrtRawFN_small_cov_write_mask; // @[Coverage map for DivSqrtRawFN_small]
  wire  DivSqrtRawFN_small_cov_write_en; // @[Coverage map for DivSqrtRawFN_small]
  reg [29:0] DivSqrtRawFN_small_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_15;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  sqrtOp_Z_shl;
  wire [4:0] sqrtOp_Z_pad;
  wire [1:0] mux_cond_0_shl;
  wire [4:0] mux_cond_0_pad;
  wire [2:0] mux_cond_1_shl;
  wire [4:0] mux_cond_1_pad;
  wire [3:0] mux_cond_2_shl;
  wire [4:0] mux_cond_2_pad;
  wire [4:0] mux_cond_3_shl;
  wire [4:0] mux_cond_3_pad;
  wire [4:0] DivSqrtRawFN_small_xor1;
  wire [4:0] DivSqrtRawFN_small_xor6;
  wire [4:0] DivSqrtRawFN_small_xor2;
  wire [4:0] DivSqrtRawFN_small_xor0;
  assign _T = io_a_isZero & io_b_isZero; // @[DivSqrtRecFN_small.scala 251:24]
  assign _T_1 = io_a_isInf & io_b_isInf; // @[DivSqrtRecFN_small.scala 251:59]
  assign notSigNaNIn_invalidExc_S_div = _T | _T_1; // @[DivSqrtRecFN_small.scala 251:42]
  assign _T_4 = ~io_a_isNaN & ~io_a_isZero; // @[DivSqrtRecFN_small.scala 253:24]
  assign notSigNaNIn_invalidExc_S_sqrt = _T_4 & io_a_sign; // @[DivSqrtRecFN_small.scala 253:43]
  assign _T_7 = io_a_isNaN & ~io_a_sig[22]; // @[common.scala 81:46]
  assign _T_8 = _T_7 | notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 256:38]
  assign _T_14 = io_b_isNaN & ~io_b_sig[22]; // @[common.scala 81:46]
  assign _T_15 = _T_7 | _T_14; // @[DivSqrtRecFN_small.scala 257:38]
  assign _T_16 = _T_15 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 257:66]
  assign _T_19 = ~io_a_isNaN & ~io_a_isInf; // @[DivSqrtRecFN_small.scala 259:33]
  assign _T_20 = _T_19 & io_b_isZero; // @[DivSqrtRecFN_small.scala 259:51]
  assign _T_21 = _T_16 | _T_20; // @[DivSqrtRecFN_small.scala 258:46]
  assign _T_22 = io_a_isNaN | notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 263:26]
  assign _T_23 = io_a_isNaN | io_b_isNaN; // @[DivSqrtRecFN_small.scala 264:26]
  assign _T_24 = _T_23 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 264:42]
  assign _T_25 = io_a_isInf | io_b_isZero; // @[DivSqrtRecFN_small.scala 266:63]
  assign _T_26 = io_a_isZero | io_b_isInf; // @[DivSqrtRecFN_small.scala 267:64]
  assign _T_28 = ~io_sqrtOp & io_b_sign; // @[DivSqrtRecFN_small.scala 268:45]
  assign sign_S = io_a_sign ^ _T_28; // @[DivSqrtRecFN_small.scala 268:30]
  assign _T_29 = io_a_isNaN | io_a_isInf; // @[DivSqrtRecFN_small.scala 270:39]
  assign specialCaseA_S = _T_29 | io_a_isZero; // @[DivSqrtRecFN_small.scala 270:55]
  assign _T_30 = io_b_isNaN | io_b_isInf; // @[DivSqrtRecFN_small.scala 271:39]
  assign specialCaseB_S = _T_30 | io_b_isZero; // @[DivSqrtRecFN_small.scala 271:55]
  assign normalCase_S_div = ~specialCaseA_S & ~specialCaseB_S; // @[DivSqrtRecFN_small.scala 272:45]
  assign normalCase_S_sqrt = ~specialCaseA_S & ~io_a_sign; // @[DivSqrtRecFN_small.scala 273:46]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[DivSqrtRecFN_small.scala 274:27]
  assign _T_39 = {io_b_sExp[8],~io_b_sExp[7:0]}; // @[DivSqrtRecFN_small.scala 278:71]
  assign _GEN_13 = {{1{_T_39[8]}},_T_39}; // @[DivSqrtRecFN_small.scala 277:21]
  assign sExpQuot_S_div = $signed(io_a_sExp) + $signed(_GEN_13); // @[DivSqrtRecFN_small.scala 277:21]
  assign _T_40 = 11'sh1c0 <= $signed(sExpQuot_S_div); // @[DivSqrtRecFN_small.scala 281:48]
  assign _T_42 = _T_40 ? 4'h6 : sExpQuot_S_div[9:6]; // @[DivSqrtRecFN_small.scala 281:16]
  assign sSatExpQuot_S_div = {_T_42,sExpQuot_S_div[5:0]}; // @[DivSqrtRecFN_small.scala 286:11]
  assign evenSqrt_S = io_sqrtOp & ~io_a_sExp[0]; // @[DivSqrtRecFN_small.scala 288:32]
  assign oddSqrt_S = io_sqrtOp & io_a_sExp[0]; // @[DivSqrtRecFN_small.scala 289:32]
  assign idle = cycleNum[0]; // @[DivSqrtRecFN_small.scala 293:24]
  assign inReady = idle | cycleNum[1]; // @[DivSqrtRecFN_small.scala 294:24]
  assign entering = inReady & io_inValid; // @[DivSqrtRecFN_small.scala 295:28]
  assign entering_normalCase = entering & normalCase_S; // @[DivSqrtRecFN_small.scala 296:40]
  assign skipCycle2 = cycleNum[3] & sigX_Z[25]; // @[DivSqrtRecFN_small.scala 298:34]
  assign _T_52 = ~idle | entering; // @[DivSqrtRecFN_small.scala 300:18]
  assign _T_54 = entering & ~normalCase_S; // @[DivSqrtRecFN_small.scala 302:26]
  assign _T_55 = _T_54 ? 2'h2 : 2'h0; // @[DivSqrtRecFN_small.scala 302:16]
  assign _T_57 = io_a_sExp[0] ? 26'h1000000 : 26'h2000000; // @[DivSqrtRecFN_small.scala 305:24]
  assign _T_58 = io_sqrtOp ? {{1'd0}, _T_57} : 27'h4000000; // @[DivSqrtRecFN_small.scala 304:20]
  assign _T_59 = entering_normalCase ? _T_58 : 27'h0; // @[DivSqrtRecFN_small.scala 303:16]
  assign _GEN_14 = {{25'd0}, _T_55}; // @[DivSqrtRecFN_small.scala 302:59]
  assign _T_60 = _GEN_14 | _T_59; // @[DivSqrtRecFN_small.scala 302:59]
  assign _T_63 = ~entering & ~skipCycle2; // @[DivSqrtRecFN_small.scala 310:28]
  assign _T_65 = _T_63 ? cycleNum[26:1] : 26'h0; // @[DivSqrtRecFN_small.scala 310:16]
  assign _GEN_15 = {{1'd0}, _T_65}; // @[DivSqrtRecFN_small.scala 309:15]
  assign _T_66 = _T_60 | _GEN_15; // @[DivSqrtRecFN_small.scala 309:15]
  assign _T_67 = skipCycle2 ? 2'h2 : 2'h0; // @[DivSqrtRecFN_small.scala 311:16]
  assign _GEN_16 = {{25'd0}, _T_67}; // @[DivSqrtRecFN_small.scala 310:63]
  assign _T_68 = _T_66 | _GEN_16; // @[DivSqrtRecFN_small.scala 310:63]
  assign _T_69 = io_a_sExp[9:1]; // @[DivSqrtRecFN_small.scala 329:29]
  assign _T_70 = $signed(_T_69) + 9'sh80; // @[DivSqrtRecFN_small.scala 329:34]
  assign _T_73 = entering_normalCase & ~io_sqrtOp; // @[DivSqrtRecFN_small.scala 334:31]
  assign _T_76 = inReady & ~oddSqrt_S; // @[DivSqrtRecFN_small.scala 341:21]
  assign _T_77 = {io_a_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 341:47]
  assign _T_78 = _T_76 ? _T_77 : 26'h0; // @[DivSqrtRecFN_small.scala 341:12]
  assign _T_79 = inReady & oddSqrt_S; // @[DivSqrtRecFN_small.scala 342:21]
  assign _T_82 = io_a_sig[23:22] - 2'h1; // @[DivSqrtRecFN_small.scala 343:56]
  assign _T_84 = {io_a_sig[21:0], 3'h0}; // @[DivSqrtRecFN_small.scala 344:44]
  assign _T_85 = {_T_82,_T_84}; // @[Cat.scala 29:58]
  assign _T_86 = _T_79 ? _T_85 : 27'h0; // @[DivSqrtRecFN_small.scala 342:12]
  assign _GEN_17 = {{1'd0}, _T_78}; // @[DivSqrtRecFN_small.scala 341:57]
  assign _T_87 = _GEN_17 | _T_86; // @[DivSqrtRecFN_small.scala 341:57]
  assign _T_89 = {rem_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 348:29]
  assign _T_90 = inReady ? 27'h0 : _T_89; // @[DivSqrtRecFN_small.scala 348:12]
  assign rem = _T_87 | _T_90; // @[DivSqrtRecFN_small.scala 347:11]
  assign bitMask = cycleNum[26:2]; // @[DivSqrtRecFN_small.scala 349:27]
  assign _T_92 = inReady & ~io_sqrtOp; // @[DivSqrtRecFN_small.scala 351:21]
  assign _T_93 = {io_b_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 351:47]
  assign _T_94 = _T_92 ? _T_93 : 26'h0; // @[DivSqrtRecFN_small.scala 351:12]
  assign _T_95 = inReady & evenSqrt_S; // @[DivSqrtRecFN_small.scala 352:21]
  assign _T_96 = _T_95 ? 25'h1000000 : 25'h0; // @[DivSqrtRecFN_small.scala 352:12]
  assign _GEN_18 = {{1'd0}, _T_96}; // @[DivSqrtRecFN_small.scala 351:73]
  assign _T_97 = _T_94 | _GEN_18; // @[DivSqrtRecFN_small.scala 351:73]
  assign _T_99 = _T_79 ? 26'h2800000 : 26'h0; // @[DivSqrtRecFN_small.scala 353:12]
  assign _T_100 = _T_97 | _T_99; // @[DivSqrtRecFN_small.scala 352:73]
  assign _T_103 = ~inReady & ~sqrtOp_Z; // @[DivSqrtRecFN_small.scala 354:23]
  assign _T_104 = {1'h1,fractB_Z}; // @[Cat.scala 29:58]
  assign _T_105 = {_T_104, 1'h0}; // @[DivSqrtRecFN_small.scala 354:56]
  assign _T_106 = _T_103 ? _T_105 : 25'h0; // @[DivSqrtRecFN_small.scala 354:12]
  assign _GEN_19 = {{1'd0}, _T_106}; // @[DivSqrtRecFN_small.scala 353:73]
  assign _T_107 = _T_100 | _GEN_19; // @[DivSqrtRecFN_small.scala 353:73]
  assign _T_109 = ~inReady & sqrtOp_Z; // @[DivSqrtRecFN_small.scala 355:23]
  assign _T_110 = {sigX_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 355:44]
  assign _GEN_20 = {{2'd0}, bitMask}; // @[DivSqrtRecFN_small.scala 355:48]
  assign _T_111 = _T_110 | _GEN_20; // @[DivSqrtRecFN_small.scala 355:48]
  assign _T_112 = _T_109 ? _T_111 : 27'h0; // @[DivSqrtRecFN_small.scala 355:12]
  assign _GEN_21 = {{1'd0}, _T_107}; // @[DivSqrtRecFN_small.scala 354:73]
  assign trialTerm = _GEN_21 | _T_112; // @[DivSqrtRecFN_small.scala 354:73]
  assign _T_113 = {1'b0,$signed(rem)}; // @[DivSqrtRecFN_small.scala 356:24]
  assign _T_114 = {1'b0,$signed(trialTerm)}; // @[DivSqrtRecFN_small.scala 356:41]
  assign trialRem = $signed(_T_113) - $signed(_T_114); // @[DivSqrtRecFN_small.scala 356:29]
  assign newBit = 28'sh0 <= $signed(trialRem); // @[DivSqrtRecFN_small.scala 357:23]
  assign _T_118 = idle | cycleNum[2]; // @[DivSqrtRecFN_small.scala 359:41]
  assign _T_120 = entering_normalCase | ~_T_118; // @[DivSqrtRecFN_small.scala 359:31]
  assign _T_121 = $signed(_T_113) - $signed(_T_114); // @[DivSqrtRecFN_small.scala 360:39]
  assign _T_122 = newBit ? _T_121 : {{1'd0}, rem}; // @[DivSqrtRecFN_small.scala 360:21]
  assign _GEN_10 = _T_120 ? _T_122 : {{2'd0}, rem_Z}; // @[DivSqrtRecFN_small.scala 359:58]
  assign _T_124 = ~inReady & newBit; // @[DivSqrtRecFN_small.scala 362:45]
  assign _T_125 = entering_normalCase | _T_124; // @[DivSqrtRecFN_small.scala 362:31]
  assign _T_126 = $signed(trialRem) != 28'sh0; // @[DivSqrtRecFN_small.scala 363:35]
  assign _T_129 = {newBit, 25'h0}; // @[DivSqrtRecFN_small.scala 365:47]
  assign _T_130 = _T_92 ? _T_129 : 26'h0; // @[DivSqrtRecFN_small.scala 365:16]
  assign _T_131 = inReady & io_sqrtOp; // @[DivSqrtRecFN_small.scala 366:25]
  assign _T_132 = _T_131 ? 25'h1000000 : 25'h0; // @[DivSqrtRecFN_small.scala 366:16]
  assign _GEN_22 = {{1'd0}, _T_132}; // @[DivSqrtRecFN_small.scala 365:71]
  assign _T_133 = _T_130 | _GEN_22; // @[DivSqrtRecFN_small.scala 365:71]
  assign _T_135 = {newBit, 23'h0}; // @[DivSqrtRecFN_small.scala 367:47]
  assign _T_136 = _T_79 ? _T_135 : 24'h0; // @[DivSqrtRecFN_small.scala 367:16]
  assign _GEN_23 = {{2'd0}, _T_136}; // @[DivSqrtRecFN_small.scala 366:71]
  assign _T_137 = _T_133 | _GEN_23; // @[DivSqrtRecFN_small.scala 366:71]
  assign _GEN_24 = {{1'd0}, bitMask}; // @[DivSqrtRecFN_small.scala 368:48]
  assign _T_139 = sigX_Z | _GEN_24; // @[DivSqrtRecFN_small.scala 368:48]
  assign _T_140 = inReady ? 26'h0 : _T_139; // @[DivSqrtRecFN_small.scala 368:16]
  assign _T_141 = _T_137 | _T_140; // @[DivSqrtRecFN_small.scala 367:71]
  assign _GEN_25 = {{26'd0}, notZeroRem_Z}; // @[DivSqrtRecFN_small.scala 385:35]
  assign io_inReady = idle | cycleNum[1]; // @[DivSqrtRecFN_small.scala 314:16]
  assign io_rawOutValid_div = cycleNum[1] & ~sqrtOp_Z; // @[DivSqrtRecFN_small.scala 375:25]
  assign io_rawOutValid_sqrt = cycleNum[1] & sqrtOp_Z; // @[DivSqrtRecFN_small.scala 376:25]
  assign io_roundingModeOut = roundingMode_Z; // @[DivSqrtRecFN_small.scala 377:25]
  assign io_invalidExc = majorExc_Z & isNaN_Z; // @[DivSqrtRecFN_small.scala 378:22]
  assign io_infiniteExc = majorExc_Z & ~isNaN_Z; // @[DivSqrtRecFN_small.scala 379:22]
  assign io_rawOut_isNaN = isNaN_Z; // @[DivSqrtRecFN_small.scala 380:22]
  assign io_rawOut_isInf = isInf_Z; // @[DivSqrtRecFN_small.scala 381:22]
  assign io_rawOut_isZero = isZero_Z; // @[DivSqrtRecFN_small.scala 382:22]
  assign io_rawOut_sign = sign_Z; // @[DivSqrtRecFN_small.scala 383:22]
  assign io_rawOut_sExp = sExp_Z; // @[DivSqrtRecFN_small.scala 384:22]
  assign io_rawOut_sig = _T_110 | _GEN_25; // @[DivSqrtRecFN_small.scala 385:22]
  assign DivSqrtRawFN_small_cov_read_addr = DivSqrtRawFN_small_state;
  assign DivSqrtRawFN_small_cov_read_data = DivSqrtRawFN_small_cov[DivSqrtRawFN_small_cov_read_addr]; // @[Coverage map for DivSqrtRawFN_small]
  assign DivSqrtRawFN_small_cov_write_data = 1'h1;
  assign DivSqrtRawFN_small_cov_write_addr = DivSqrtRawFN_small_state;
  assign DivSqrtRawFN_small_cov_write_mask = 1'h1;
  assign DivSqrtRawFN_small_cov_write_en = 1'h1;
  assign mux_cond_0 = _T_125;
  assign mux_cond_1 = newBit;
  assign mux_cond_2 = _T_63;
  assign mux_cond_3 = skipCycle2;
  assign sqrtOp_Z_shl = sqrtOp_Z;
  assign sqrtOp_Z_pad = {4'h0,sqrtOp_Z_shl};
  assign mux_cond_0_shl = {mux_cond_0, 1'h0};
  assign mux_cond_0_pad = {3'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 2'h0};
  assign mux_cond_1_pad = {2'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 3'h0};
  assign mux_cond_2_pad = {1'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 4'h0};
  assign mux_cond_3_pad = mux_cond_3_shl;
  assign DivSqrtRawFN_small_xor1 = sqrtOp_Z_pad ^ mux_cond_0_pad;
  assign DivSqrtRawFN_small_xor6 = mux_cond_2_pad ^ mux_cond_3_pad;
  assign DivSqrtRawFN_small_xor2 = mux_cond_1_pad ^ DivSqrtRawFN_small_xor6;
  assign DivSqrtRawFN_small_xor0 = DivSqrtRawFN_small_xor1 ^ DivSqrtRawFN_small_xor2;
  assign io_covSum = DivSqrtRawFN_small_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  majorExc_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isNaN_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  isInf_Z = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  isZero_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sign_Z = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sExp_Z = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  fractB_Z = _RAND_8[22:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  roundingMode_Z = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  rem_Z = _RAND_10[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  notZeroRem_Z = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  sigX_Z = _RAND_12[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  DivSqrtRawFN_small_state = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    DivSqrtRawFN_small_cov[initvar] = _RAND_14[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  DivSqrtRawFN_small_covSum = _RAND_15[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      cycleNum <= 27'h0;
    end else if (reset) begin
      cycleNum <= 27'h1;
    end else if (_T_52) begin
      cycleNum <= _T_68;
    end
    if (metaReset) begin
      sqrtOp_Z <= 1'h0;
    end else if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (metaReset) begin
      majorExc_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        majorExc_Z <= _T_8;
      end else begin
        majorExc_Z <= _T_21;
      end
    end
    if (metaReset) begin
      isNaN_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isNaN_Z <= _T_22;
      end else begin
        isNaN_Z <= _T_24;
      end
    end
    if (metaReset) begin
      isInf_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isInf_Z <= io_a_isInf;
      end else begin
        isInf_Z <= _T_25;
      end
    end
    if (metaReset) begin
      isZero_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= io_a_isZero;
      end else begin
        isZero_Z <= _T_26;
      end
    end
    if (metaReset) begin
      sign_Z <= 1'h0;
    end else if (entering) begin
      sign_Z <= sign_S;
    end
    if (metaReset) begin
      sExp_Z <= 10'h0;
    end else if (entering_normalCase) begin
      if (io_sqrtOp) begin
        sExp_Z <= _T_70;
      end else begin
        sExp_Z <= sSatExpQuot_S_div;
      end
    end
    if (metaReset) begin
      fractB_Z <= 23'h0;
    end else if (_T_73) begin
      fractB_Z <= io_b_sig[22:0];
    end
    if (metaReset) begin
      roundingMode_Z <= 3'h0;
    end else if (entering_normalCase) begin
      roundingMode_Z <= io_roundingMode;
    end
    if (metaReset) begin
      rem_Z <= 26'h0;
    end else begin
      rem_Z <= _GEN_10[25:0];
    end
    if (metaReset) begin
      notZeroRem_Z <= 1'h0;
    end else if (_T_125) begin
      notZeroRem_Z <= _T_126;
    end
    if (metaReset) begin
      sigX_Z <= 26'h0;
    end else if (_T_125) begin
      sigX_Z <= _T_141;
    end
    DivSqrtRawFN_small_state <= DivSqrtRawFN_small_xor0;
    if (!(DivSqrtRawFN_small_cov_read_data)) begin
      DivSqrtRawFN_small_covSum <= DivSqrtRawFN_small_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(DivSqrtRawFN_small_cov_write_en & DivSqrtRawFN_small_cov_write_mask) begin
      DivSqrtRawFN_small_cov[DivSqrtRawFN_small_cov_write_addr] <= DivSqrtRawFN_small_cov_write_data; // @[Coverage map for DivSqrtRawFN_small]
    end
  end
endmodule
module RoundAnyRawFNToRecFN_5(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire  doShiftSigDown1; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire  _T_5; // @[primitives.scala 57:25]
  wire  _T_7; // @[primitives.scala 57:25]
  wire  _T_9; // @[primitives.scala 57:25]
  wire [5:0] _T_10; // @[primitives.scala 58:26]
  wire [64:0] _T_11; // @[primitives.scala 77:58]
  wire [15:0] _T_17; // @[Bitwise.scala 103:31]
  wire [15:0] _T_19; // @[Bitwise.scala 103:65]
  wire [15:0] _T_21; // @[Bitwise.scala 103:75]
  wire [15:0] _T_22; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_0; // @[Bitwise.scala 103:31]
  wire [15:0] _T_27; // @[Bitwise.scala 103:31]
  wire [15:0] _T_29; // @[Bitwise.scala 103:65]
  wire [15:0] _T_31; // @[Bitwise.scala 103:75]
  wire [15:0] _T_32; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [15:0] _T_37; // @[Bitwise.scala 103:31]
  wire [15:0] _T_39; // @[Bitwise.scala 103:65]
  wire [15:0] _T_41; // @[Bitwise.scala 103:75]
  wire [15:0] _T_42; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [15:0] _T_47; // @[Bitwise.scala 103:31]
  wire [15:0] _T_49; // @[Bitwise.scala 103:65]
  wire [15:0] _T_51; // @[Bitwise.scala 103:75]
  wire [15:0] _T_52; // @[Bitwise.scala 103:39]
  wire [21:0] _T_69; // @[Cat.scala 29:58]
  wire [21:0] _T_71; // @[primitives.scala 74:21]
  wire [24:0] _T_73; // @[Cat.scala 29:58]
  wire [2:0] _T_83; // @[Cat.scala 29:58]
  wire [2:0] _T_84; // @[primitives.scala 61:24]
  wire [24:0] _T_85; // @[primitives.scala 66:24]
  wire [24:0] _T_86; // @[primitives.scala 61:24]
  wire [24:0] _GEN_3; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [24:0] _T_87; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [26:0] _T_88; // @[Cat.scala 29:58]
  wire [26:0] _T_90; // @[Cat.scala 29:58]
  wire [26:0] _T_92; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [26:0] _T_93; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_94; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _T_95; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_96; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  _T_97; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_98; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_99; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_100; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_101; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [26:0] _T_102; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _T_104; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_105; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_107; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [25:0] _T_109; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _T_111; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _T_113; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_115; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [25:0] _T_117; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [25:0] _GEN_4; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_118; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_119; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_121; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [9:0] _GEN_5; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [10:0] _T_122; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _T_127; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  _T_132; // @[RoundAnyRawFNToRecFN.scala 201:16]
  wire  _T_134; // @[RoundAnyRawFNToRecFN.scala 203:30]
  wire  _T_136; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _T_137; // @[RoundAnyRawFNToRecFN.scala 203:49]
  wire  _T_139; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _T_140; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  _T_141; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire  _T_144; // @[RoundAnyRawFNToRecFN.scala 209:16]
  wire [1:0] _T_145; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _T_146; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _T_147; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _T_150; // @[RoundAnyRawFNToRecFN.scala 219:30]
  wire  _T_151; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _T_155; // @[RoundAnyRawFNToRecFN.scala 221:39]
  wire  _T_157; // @[RoundAnyRawFNToRecFN.scala 220:77]
  wire  _T_158; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _T_159; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _T_160; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _T_162; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 234:49]
  wire  _T_167; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _T_169; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _T_171; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _T_172; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _T_174; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _T_175; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [8:0] _T_176; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] _T_178; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [8:0] _T_180; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [8:0] _T_182; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [8:0] _T_183; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [8:0] _T_185; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [8:0] _T_186; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [8:0] _T_188; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [8:0] _T_189; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [8:0] _T_190; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [8:0] _T_191; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [8:0] _T_192; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [8:0] _T_193; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [8:0] _T_194; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [8:0] _T_195; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_196; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _T_197; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [22:0] _T_198; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [22:0] _T_199; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [22:0] _T_201; // @[Bitwise.scala 72:12]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [9:0] _T_202; // @[Cat.scala 29:58]
  wire [1:0] _T_204; // @[Cat.scala 29:58]
  wire [2:0] _T_206; // @[Cat.scala 29:58]
  wire [29:0] RoundAnyRawFNToRecFN_5_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign doShiftSigDown1 = io_in_sig[26]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  assign _T_5 = ~io_in_sExp[8]; // @[primitives.scala 57:25]
  assign _T_7 = ~io_in_sExp[7]; // @[primitives.scala 57:25]
  assign _T_9 = ~io_in_sExp[6]; // @[primitives.scala 57:25]
  assign _T_10 = ~io_in_sExp[5:0]; // @[primitives.scala 58:26]
  assign _T_11 = -65'sh10000000000000000 >>> _T_10; // @[primitives.scala 77:58]
  assign _T_17 = {{8'd0}, _T_11[57:50]}; // @[Bitwise.scala 103:31]
  assign _T_19 = {_T_11[49:42], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_21 = _T_19 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_22 = _T_17 | _T_21; // @[Bitwise.scala 103:39]
  assign _GEN_0 = {{4'd0}, _T_22[15:4]}; // @[Bitwise.scala 103:31]
  assign _T_27 = _GEN_0 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_29 = {_T_22[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_31 = _T_29 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_32 = _T_27 | _T_31; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{2'd0}, _T_32[15:2]}; // @[Bitwise.scala 103:31]
  assign _T_37 = _GEN_1 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_39 = {_T_32[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_41 = _T_39 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_42 = _T_37 | _T_41; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{1'd0}, _T_42[15:1]}; // @[Bitwise.scala 103:31]
  assign _T_47 = _GEN_2 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_49 = {_T_42[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_51 = _T_49 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_52 = _T_47 | _T_51; // @[Bitwise.scala 103:39]
  assign _T_69 = {_T_52,_T_11[58],_T_11[59],_T_11[60],_T_11[61],_T_11[62],_T_11[63]}; // @[Cat.scala 29:58]
  assign _T_71 = _T_9 ? 22'h0 : ~_T_69; // @[primitives.scala 74:21]
  assign _T_73 = {~_T_71,3'h7}; // @[Cat.scala 29:58]
  assign _T_83 = {_T_11[0],_T_11[1],_T_11[2]}; // @[Cat.scala 29:58]
  assign _T_84 = _T_9 ? _T_83 : 3'h0; // @[primitives.scala 61:24]
  assign _T_85 = _T_7 ? _T_73 : {{22'd0}, _T_84}; // @[primitives.scala 66:24]
  assign _T_86 = _T_5 ? _T_85 : 25'h0; // @[primitives.scala 61:24]
  assign _GEN_3 = {{24'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_87 = _T_86 | _GEN_3; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_88 = {_T_87,2'h3}; // @[Cat.scala 29:58]
  assign _T_90 = {1'h0,_T_88[26:1]}; // @[Cat.scala 29:58]
  assign _T_92 = ~_T_90 & _T_88; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _T_93 = io_in_sig & _T_92; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_94 = |_T_93; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_95 = io_in_sig & _T_90; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_96 = |_T_95; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign _T_97 = _T_94 | _T_96; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_98 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_99 = _T_98 & _T_94; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_100 = roundMagUp & _T_97; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_101 = _T_99 | _T_100; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_102 = io_in_sig | _T_88; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_104 = _T_102[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_105 = roundingMode_near_even & _T_94; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_107 = _T_105 & ~_T_96; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_109 = _T_107 ? _T_88[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_111 = _T_104 & ~_T_109; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_113 = io_in_sig & ~_T_88; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_115 = roundingMode_odd & _T_97; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_117 = _T_115 ? _T_92[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_4 = {{1'd0}, _T_113[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_118 = _GEN_4 | _T_117; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_119 = _T_101 ? _T_111 : _T_118; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_121 = {1'b0,$signed(_T_119[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_5 = {{7{_T_121[2]}},_T_121}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_122 = $signed(io_in_sExp) + $signed(_GEN_5); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_122[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = doShiftSigDown1 ? _T_119[23:1] : _T_119[22:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  assign _T_127 = _T_122[10:7]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_T_127) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(_T_122) < 11'sh6b; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign _T_132 = doShiftSigDown1 ? io_in_sig[2] : io_in_sig[1]; // @[RoundAnyRawFNToRecFN.scala 201:16]
  assign _T_134 = doShiftSigDown1 & io_in_sig[2]; // @[RoundAnyRawFNToRecFN.scala 203:30]
  assign _T_136 = |io_in_sig[1:0]; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign _T_137 = _T_134 | _T_136; // @[RoundAnyRawFNToRecFN.scala 203:49]
  assign _T_139 = _T_98 & _T_132; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _T_140 = roundMagUp & _T_137; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign _T_141 = _T_139 | _T_140; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign _T_144 = doShiftSigDown1 ? _T_119[25] : _T_119[24]; // @[RoundAnyRawFNToRecFN.scala 209:16]
  assign _T_145 = io_in_sExp[9:8]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _T_146 = $signed(_T_145) <= 2'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _T_147 = _T_97 & _T_146; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _T_150 = doShiftSigDown1 ? _T_88[3] : _T_88[2]; // @[RoundAnyRawFNToRecFN.scala 219:30]
  assign _T_151 = _T_147 & _T_150; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _T_155 = doShiftSigDown1 ? _T_88[4] : _T_88[3]; // @[RoundAnyRawFNToRecFN.scala 221:39]
  assign _T_157 = io_detectTininess & ~_T_155; // @[RoundAnyRawFNToRecFN.scala 220:77]
  assign _T_158 = _T_157 & _T_144; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _T_159 = _T_158 & _T_94; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _T_160 = _T_159 & _T_141; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _T_162 = _T_151 & ~_T_160; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _T_162; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | _T_97; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 234:49]
  assign _T_167 = ~isNaNOut & ~notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _T_167 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _T_169 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _T_169; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _T_98 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _T_171 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _T_172 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _T_171 & _T_172; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _T_174 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | _T_174; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _T_175 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _T_176 = _T_175 ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_178 = common_expOut & ~_T_176; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_180 = pegMinNonzeroMagOut ? 9'h194 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _T_182 = _T_178 & ~_T_180; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _T_183 = pegMaxFiniteMagOut ? 9'h80 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _T_185 = _T_182 & ~_T_183; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _T_186 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_188 = _T_185 & ~_T_186; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_189 = pegMinNonzeroMagOut ? 9'h6b : 9'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _T_190 = _T_188 | _T_189; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _T_191 = pegMaxFiniteMagOut ? 9'h17f : 9'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _T_192 = _T_190 | _T_191; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _T_193 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _T_194 = _T_192 | _T_193; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_195 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _T_194 | _T_195; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _T_196 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _T_197 = _T_196 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _T_198 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _T_199 = _T_197 ? _T_198 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_201 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0; // @[Bitwise.scala 72:12]
  assign fractOut = _T_199 | _T_201; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign _T_202 = {signOut,expOut}; // @[Cat.scala 29:58]
  assign _T_204 = {underflow,inexact}; // @[Cat.scala 29:58]
  assign _T_206 = {io_invalidExc,io_infiniteExc,overflow}; // @[Cat.scala 29:58]
  assign io_out = {_T_202,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_206,_T_204}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_5_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_5_covSum;
  assign metaAssert = 1'h0;
endmodule
module DivSqrtRawFN_small_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [12:0] io_a_sExp,
  input  [53:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [12:0] io_b_sExp,
  input  [53:0] io_b_sig,
  input  [2:0]  io_roundingMode,
  output        io_rawOutValid_div,
  output        io_rawOutValid_sqrt,
  output [2:0]  io_roundingModeOut,
  output        io_invalidExc,
  output        io_infiniteExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [12:0] io_rawOut_sExp,
  output [55:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [55:0] cycleNum; // @[DivSqrtRecFN_small.scala 223:33]
  reg [63:0] _RAND_0;
  reg  sqrtOp_Z; // @[DivSqrtRecFN_small.scala 225:29]
  reg [31:0] _RAND_1;
  reg  majorExc_Z; // @[DivSqrtRecFN_small.scala 226:29]
  reg [31:0] _RAND_2;
  reg  isNaN_Z; // @[DivSqrtRecFN_small.scala 228:29]
  reg [31:0] _RAND_3;
  reg  isInf_Z; // @[DivSqrtRecFN_small.scala 229:29]
  reg [31:0] _RAND_4;
  reg  isZero_Z; // @[DivSqrtRecFN_small.scala 230:29]
  reg [31:0] _RAND_5;
  reg  sign_Z; // @[DivSqrtRecFN_small.scala 231:29]
  reg [31:0] _RAND_6;
  reg [12:0] sExp_Z; // @[DivSqrtRecFN_small.scala 232:29]
  reg [31:0] _RAND_7;
  reg [51:0] fractB_Z; // @[DivSqrtRecFN_small.scala 233:29]
  reg [63:0] _RAND_8;
  reg [2:0] roundingMode_Z; // @[DivSqrtRecFN_small.scala 234:29]
  reg [31:0] _RAND_9;
  reg [54:0] rem_Z; // @[DivSqrtRecFN_small.scala 240:29]
  reg [63:0] _RAND_10;
  reg  notZeroRem_Z; // @[DivSqrtRecFN_small.scala 241:29]
  reg [31:0] _RAND_11;
  reg [54:0] sigX_Z; // @[DivSqrtRecFN_small.scala 242:29]
  reg [63:0] _RAND_12;
  wire  _T; // @[DivSqrtRecFN_small.scala 251:24]
  wire  _T_1; // @[DivSqrtRecFN_small.scala 251:59]
  wire  notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 251:42]
  wire  _T_4; // @[DivSqrtRecFN_small.scala 253:24]
  wire  notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 253:43]
  wire  _T_7; // @[common.scala 81:46]
  wire  _T_8; // @[DivSqrtRecFN_small.scala 256:38]
  wire  _T_14; // @[common.scala 81:46]
  wire  _T_15; // @[DivSqrtRecFN_small.scala 257:38]
  wire  _T_16; // @[DivSqrtRecFN_small.scala 257:66]
  wire  _T_19; // @[DivSqrtRecFN_small.scala 259:33]
  wire  _T_20; // @[DivSqrtRecFN_small.scala 259:51]
  wire  _T_21; // @[DivSqrtRecFN_small.scala 258:46]
  wire  _T_22; // @[DivSqrtRecFN_small.scala 263:26]
  wire  _T_23; // @[DivSqrtRecFN_small.scala 264:26]
  wire  _T_24; // @[DivSqrtRecFN_small.scala 264:42]
  wire  _T_25; // @[DivSqrtRecFN_small.scala 266:63]
  wire  _T_26; // @[DivSqrtRecFN_small.scala 267:64]
  wire  _T_28; // @[DivSqrtRecFN_small.scala 268:45]
  wire  sign_S; // @[DivSqrtRecFN_small.scala 268:30]
  wire  _T_29; // @[DivSqrtRecFN_small.scala 270:39]
  wire  specialCaseA_S; // @[DivSqrtRecFN_small.scala 270:55]
  wire  _T_30; // @[DivSqrtRecFN_small.scala 271:39]
  wire  specialCaseB_S; // @[DivSqrtRecFN_small.scala 271:55]
  wire  normalCase_S_div; // @[DivSqrtRecFN_small.scala 272:45]
  wire  normalCase_S_sqrt; // @[DivSqrtRecFN_small.scala 273:46]
  wire  normalCase_S; // @[DivSqrtRecFN_small.scala 274:27]
  wire [11:0] _T_39; // @[DivSqrtRecFN_small.scala 278:71]
  wire [12:0] _GEN_13; // @[DivSqrtRecFN_small.scala 277:21]
  wire [13:0] sExpQuot_S_div; // @[DivSqrtRecFN_small.scala 277:21]
  wire  _T_40; // @[DivSqrtRecFN_small.scala 281:48]
  wire [3:0] _T_42; // @[DivSqrtRecFN_small.scala 281:16]
  wire [12:0] sSatExpQuot_S_div; // @[DivSqrtRecFN_small.scala 286:11]
  wire  evenSqrt_S; // @[DivSqrtRecFN_small.scala 288:32]
  wire  oddSqrt_S; // @[DivSqrtRecFN_small.scala 289:32]
  wire  idle; // @[DivSqrtRecFN_small.scala 293:24]
  wire  inReady; // @[DivSqrtRecFN_small.scala 294:24]
  wire  entering; // @[DivSqrtRecFN_small.scala 295:28]
  wire  entering_normalCase; // @[DivSqrtRecFN_small.scala 296:40]
  wire  skipCycle2; // @[DivSqrtRecFN_small.scala 298:34]
  wire  _T_52; // @[DivSqrtRecFN_small.scala 300:18]
  wire  _T_54; // @[DivSqrtRecFN_small.scala 302:26]
  wire [1:0] _T_55; // @[DivSqrtRecFN_small.scala 302:16]
  wire [54:0] _T_57; // @[DivSqrtRecFN_small.scala 305:24]
  wire [55:0] _T_58; // @[DivSqrtRecFN_small.scala 304:20]
  wire [55:0] _T_59; // @[DivSqrtRecFN_small.scala 303:16]
  wire [55:0] _GEN_14; // @[DivSqrtRecFN_small.scala 302:59]
  wire [55:0] _T_60; // @[DivSqrtRecFN_small.scala 302:59]
  wire  _T_63; // @[DivSqrtRecFN_small.scala 310:28]
  wire [54:0] _T_65; // @[DivSqrtRecFN_small.scala 310:16]
  wire [55:0] _GEN_15; // @[DivSqrtRecFN_small.scala 309:15]
  wire [55:0] _T_66; // @[DivSqrtRecFN_small.scala 309:15]
  wire [1:0] _T_67; // @[DivSqrtRecFN_small.scala 311:16]
  wire [55:0] _GEN_16; // @[DivSqrtRecFN_small.scala 310:63]
  wire [55:0] _T_68; // @[DivSqrtRecFN_small.scala 310:63]
  wire [11:0] _T_69; // @[DivSqrtRecFN_small.scala 329:29]
  wire [12:0] _T_70; // @[DivSqrtRecFN_small.scala 329:34]
  wire  _T_73; // @[DivSqrtRecFN_small.scala 334:31]
  wire  _T_76; // @[DivSqrtRecFN_small.scala 341:21]
  wire [54:0] _T_77; // @[DivSqrtRecFN_small.scala 341:47]
  wire [54:0] _T_78; // @[DivSqrtRecFN_small.scala 341:12]
  wire  _T_79; // @[DivSqrtRecFN_small.scala 342:21]
  wire [1:0] _T_82; // @[DivSqrtRecFN_small.scala 343:56]
  wire [53:0] _T_84; // @[DivSqrtRecFN_small.scala 344:44]
  wire [55:0] _T_85; // @[Cat.scala 29:58]
  wire [55:0] _T_86; // @[DivSqrtRecFN_small.scala 342:12]
  wire [55:0] _GEN_17; // @[DivSqrtRecFN_small.scala 341:57]
  wire [55:0] _T_87; // @[DivSqrtRecFN_small.scala 341:57]
  wire [55:0] _T_89; // @[DivSqrtRecFN_small.scala 348:29]
  wire [55:0] _T_90; // @[DivSqrtRecFN_small.scala 348:12]
  wire [55:0] rem; // @[DivSqrtRecFN_small.scala 347:11]
  wire [53:0] bitMask; // @[DivSqrtRecFN_small.scala 349:27]
  wire  _T_92; // @[DivSqrtRecFN_small.scala 351:21]
  wire [54:0] _T_93; // @[DivSqrtRecFN_small.scala 351:47]
  wire [54:0] _T_94; // @[DivSqrtRecFN_small.scala 351:12]
  wire  _T_95; // @[DivSqrtRecFN_small.scala 352:21]
  wire [53:0] _T_96; // @[DivSqrtRecFN_small.scala 352:12]
  wire [54:0] _GEN_18; // @[DivSqrtRecFN_small.scala 351:73]
  wire [54:0] _T_97; // @[DivSqrtRecFN_small.scala 351:73]
  wire [54:0] _T_99; // @[DivSqrtRecFN_small.scala 353:12]
  wire [54:0] _T_100; // @[DivSqrtRecFN_small.scala 352:73]
  wire  _T_103; // @[DivSqrtRecFN_small.scala 354:23]
  wire [52:0] _T_104; // @[Cat.scala 29:58]
  wire [53:0] _T_105; // @[DivSqrtRecFN_small.scala 354:56]
  wire [53:0] _T_106; // @[DivSqrtRecFN_small.scala 354:12]
  wire [54:0] _GEN_19; // @[DivSqrtRecFN_small.scala 353:73]
  wire [54:0] _T_107; // @[DivSqrtRecFN_small.scala 353:73]
  wire  _T_109; // @[DivSqrtRecFN_small.scala 355:23]
  wire [55:0] _T_110; // @[DivSqrtRecFN_small.scala 355:44]
  wire [55:0] _GEN_20; // @[DivSqrtRecFN_small.scala 355:48]
  wire [55:0] _T_111; // @[DivSqrtRecFN_small.scala 355:48]
  wire [55:0] _T_112; // @[DivSqrtRecFN_small.scala 355:12]
  wire [55:0] _GEN_21; // @[DivSqrtRecFN_small.scala 354:73]
  wire [55:0] trialTerm; // @[DivSqrtRecFN_small.scala 354:73]
  wire [56:0] _T_113; // @[DivSqrtRecFN_small.scala 356:24]
  wire [56:0] _T_114; // @[DivSqrtRecFN_small.scala 356:41]
  wire [56:0] trialRem; // @[DivSqrtRecFN_small.scala 356:29]
  wire  newBit; // @[DivSqrtRecFN_small.scala 357:23]
  wire  _T_118; // @[DivSqrtRecFN_small.scala 359:41]
  wire  _T_120; // @[DivSqrtRecFN_small.scala 359:31]
  wire [56:0] _T_121; // @[DivSqrtRecFN_small.scala 360:39]
  wire [56:0] _T_122; // @[DivSqrtRecFN_small.scala 360:21]
  wire [56:0] _GEN_10; // @[DivSqrtRecFN_small.scala 359:58]
  wire  _T_124; // @[DivSqrtRecFN_small.scala 362:45]
  wire  _T_125; // @[DivSqrtRecFN_small.scala 362:31]
  wire  _T_126; // @[DivSqrtRecFN_small.scala 363:35]
  wire [54:0] _T_129; // @[DivSqrtRecFN_small.scala 365:47]
  wire [54:0] _T_130; // @[DivSqrtRecFN_small.scala 365:16]
  wire  _T_131; // @[DivSqrtRecFN_small.scala 366:25]
  wire [53:0] _T_132; // @[DivSqrtRecFN_small.scala 366:16]
  wire [54:0] _GEN_22; // @[DivSqrtRecFN_small.scala 365:71]
  wire [54:0] _T_133; // @[DivSqrtRecFN_small.scala 365:71]
  wire [52:0] _T_135; // @[DivSqrtRecFN_small.scala 367:47]
  wire [52:0] _T_136; // @[DivSqrtRecFN_small.scala 367:16]
  wire [54:0] _GEN_23; // @[DivSqrtRecFN_small.scala 366:71]
  wire [54:0] _T_137; // @[DivSqrtRecFN_small.scala 366:71]
  wire [54:0] _GEN_24; // @[DivSqrtRecFN_small.scala 368:48]
  wire [54:0] _T_139; // @[DivSqrtRecFN_small.scala 368:48]
  wire [54:0] _T_140; // @[DivSqrtRecFN_small.scala 368:16]
  wire [54:0] _T_141; // @[DivSqrtRecFN_small.scala 367:71]
  wire [55:0] _GEN_25; // @[DivSqrtRecFN_small.scala 385:35]
  reg [4:0] DivSqrtRawFN_small_1_state; // @[Register tracking DivSqrtRawFN_small_1 state]
  reg [31:0] _RAND_13;
  reg  DivSqrtRawFN_small_1_cov [0:31]; // @[Coverage map for DivSqrtRawFN_small_1]
  reg [31:0] _RAND_14;
  wire  DivSqrtRawFN_small_1_cov_read_data; // @[Coverage map for DivSqrtRawFN_small_1]
  wire [4:0] DivSqrtRawFN_small_1_cov_read_addr; // @[Coverage map for DivSqrtRawFN_small_1]
  wire  DivSqrtRawFN_small_1_cov_write_data; // @[Coverage map for DivSqrtRawFN_small_1]
  wire [4:0] DivSqrtRawFN_small_1_cov_write_addr; // @[Coverage map for DivSqrtRawFN_small_1]
  wire  DivSqrtRawFN_small_1_cov_write_mask; // @[Coverage map for DivSqrtRawFN_small_1]
  wire  DivSqrtRawFN_small_1_cov_write_en; // @[Coverage map for DivSqrtRawFN_small_1]
  reg [29:0] DivSqrtRawFN_small_1_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_15;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  sqrtOp_Z_shl;
  wire [4:0] sqrtOp_Z_pad;
  wire [1:0] mux_cond_0_shl;
  wire [4:0] mux_cond_0_pad;
  wire [2:0] mux_cond_1_shl;
  wire [4:0] mux_cond_1_pad;
  wire [3:0] mux_cond_2_shl;
  wire [4:0] mux_cond_2_pad;
  wire [4:0] mux_cond_3_shl;
  wire [4:0] mux_cond_3_pad;
  wire [4:0] DivSqrtRawFN_small_1_xor1;
  wire [4:0] DivSqrtRawFN_small_1_xor6;
  wire [4:0] DivSqrtRawFN_small_1_xor2;
  wire [4:0] DivSqrtRawFN_small_1_xor0;
  assign _T = io_a_isZero & io_b_isZero; // @[DivSqrtRecFN_small.scala 251:24]
  assign _T_1 = io_a_isInf & io_b_isInf; // @[DivSqrtRecFN_small.scala 251:59]
  assign notSigNaNIn_invalidExc_S_div = _T | _T_1; // @[DivSqrtRecFN_small.scala 251:42]
  assign _T_4 = ~io_a_isNaN & ~io_a_isZero; // @[DivSqrtRecFN_small.scala 253:24]
  assign notSigNaNIn_invalidExc_S_sqrt = _T_4 & io_a_sign; // @[DivSqrtRecFN_small.scala 253:43]
  assign _T_7 = io_a_isNaN & ~io_a_sig[51]; // @[common.scala 81:46]
  assign _T_8 = _T_7 | notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 256:38]
  assign _T_14 = io_b_isNaN & ~io_b_sig[51]; // @[common.scala 81:46]
  assign _T_15 = _T_7 | _T_14; // @[DivSqrtRecFN_small.scala 257:38]
  assign _T_16 = _T_15 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 257:66]
  assign _T_19 = ~io_a_isNaN & ~io_a_isInf; // @[DivSqrtRecFN_small.scala 259:33]
  assign _T_20 = _T_19 & io_b_isZero; // @[DivSqrtRecFN_small.scala 259:51]
  assign _T_21 = _T_16 | _T_20; // @[DivSqrtRecFN_small.scala 258:46]
  assign _T_22 = io_a_isNaN | notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 263:26]
  assign _T_23 = io_a_isNaN | io_b_isNaN; // @[DivSqrtRecFN_small.scala 264:26]
  assign _T_24 = _T_23 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 264:42]
  assign _T_25 = io_a_isInf | io_b_isZero; // @[DivSqrtRecFN_small.scala 266:63]
  assign _T_26 = io_a_isZero | io_b_isInf; // @[DivSqrtRecFN_small.scala 267:64]
  assign _T_28 = ~io_sqrtOp & io_b_sign; // @[DivSqrtRecFN_small.scala 268:45]
  assign sign_S = io_a_sign ^ _T_28; // @[DivSqrtRecFN_small.scala 268:30]
  assign _T_29 = io_a_isNaN | io_a_isInf; // @[DivSqrtRecFN_small.scala 270:39]
  assign specialCaseA_S = _T_29 | io_a_isZero; // @[DivSqrtRecFN_small.scala 270:55]
  assign _T_30 = io_b_isNaN | io_b_isInf; // @[DivSqrtRecFN_small.scala 271:39]
  assign specialCaseB_S = _T_30 | io_b_isZero; // @[DivSqrtRecFN_small.scala 271:55]
  assign normalCase_S_div = ~specialCaseA_S & ~specialCaseB_S; // @[DivSqrtRecFN_small.scala 272:45]
  assign normalCase_S_sqrt = ~specialCaseA_S & ~io_a_sign; // @[DivSqrtRecFN_small.scala 273:46]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[DivSqrtRecFN_small.scala 274:27]
  assign _T_39 = {io_b_sExp[11],~io_b_sExp[10:0]}; // @[DivSqrtRecFN_small.scala 278:71]
  assign _GEN_13 = {{1{_T_39[11]}},_T_39}; // @[DivSqrtRecFN_small.scala 277:21]
  assign sExpQuot_S_div = $signed(io_a_sExp) + $signed(_GEN_13); // @[DivSqrtRecFN_small.scala 277:21]
  assign _T_40 = 14'she00 <= $signed(sExpQuot_S_div); // @[DivSqrtRecFN_small.scala 281:48]
  assign _T_42 = _T_40 ? 4'h6 : sExpQuot_S_div[12:9]; // @[DivSqrtRecFN_small.scala 281:16]
  assign sSatExpQuot_S_div = {_T_42,sExpQuot_S_div[8:0]}; // @[DivSqrtRecFN_small.scala 286:11]
  assign evenSqrt_S = io_sqrtOp & ~io_a_sExp[0]; // @[DivSqrtRecFN_small.scala 288:32]
  assign oddSqrt_S = io_sqrtOp & io_a_sExp[0]; // @[DivSqrtRecFN_small.scala 289:32]
  assign idle = cycleNum[0]; // @[DivSqrtRecFN_small.scala 293:24]
  assign inReady = idle | cycleNum[1]; // @[DivSqrtRecFN_small.scala 294:24]
  assign entering = inReady & io_inValid; // @[DivSqrtRecFN_small.scala 295:28]
  assign entering_normalCase = entering & normalCase_S; // @[DivSqrtRecFN_small.scala 296:40]
  assign skipCycle2 = cycleNum[3] & sigX_Z[54]; // @[DivSqrtRecFN_small.scala 298:34]
  assign _T_52 = ~idle | entering; // @[DivSqrtRecFN_small.scala 300:18]
  assign _T_54 = entering & ~normalCase_S; // @[DivSqrtRecFN_small.scala 302:26]
  assign _T_55 = _T_54 ? 2'h2 : 2'h0; // @[DivSqrtRecFN_small.scala 302:16]
  assign _T_57 = io_a_sExp[0] ? 55'h20000000000000 : 55'h40000000000000; // @[DivSqrtRecFN_small.scala 305:24]
  assign _T_58 = io_sqrtOp ? {{1'd0}, _T_57} : 56'h80000000000000; // @[DivSqrtRecFN_small.scala 304:20]
  assign _T_59 = entering_normalCase ? _T_58 : 56'h0; // @[DivSqrtRecFN_small.scala 303:16]
  assign _GEN_14 = {{54'd0}, _T_55}; // @[DivSqrtRecFN_small.scala 302:59]
  assign _T_60 = _GEN_14 | _T_59; // @[DivSqrtRecFN_small.scala 302:59]
  assign _T_63 = ~entering & ~skipCycle2; // @[DivSqrtRecFN_small.scala 310:28]
  assign _T_65 = _T_63 ? cycleNum[55:1] : 55'h0; // @[DivSqrtRecFN_small.scala 310:16]
  assign _GEN_15 = {{1'd0}, _T_65}; // @[DivSqrtRecFN_small.scala 309:15]
  assign _T_66 = _T_60 | _GEN_15; // @[DivSqrtRecFN_small.scala 309:15]
  assign _T_67 = skipCycle2 ? 2'h2 : 2'h0; // @[DivSqrtRecFN_small.scala 311:16]
  assign _GEN_16 = {{54'd0}, _T_67}; // @[DivSqrtRecFN_small.scala 310:63]
  assign _T_68 = _T_66 | _GEN_16; // @[DivSqrtRecFN_small.scala 310:63]
  assign _T_69 = io_a_sExp[12:1]; // @[DivSqrtRecFN_small.scala 329:29]
  assign _T_70 = $signed(_T_69) + 12'sh400; // @[DivSqrtRecFN_small.scala 329:34]
  assign _T_73 = entering_normalCase & ~io_sqrtOp; // @[DivSqrtRecFN_small.scala 334:31]
  assign _T_76 = inReady & ~oddSqrt_S; // @[DivSqrtRecFN_small.scala 341:21]
  assign _T_77 = {io_a_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 341:47]
  assign _T_78 = _T_76 ? _T_77 : 55'h0; // @[DivSqrtRecFN_small.scala 341:12]
  assign _T_79 = inReady & oddSqrt_S; // @[DivSqrtRecFN_small.scala 342:21]
  assign _T_82 = io_a_sig[52:51] - 2'h1; // @[DivSqrtRecFN_small.scala 343:56]
  assign _T_84 = {io_a_sig[50:0], 3'h0}; // @[DivSqrtRecFN_small.scala 344:44]
  assign _T_85 = {_T_82,_T_84}; // @[Cat.scala 29:58]
  assign _T_86 = _T_79 ? _T_85 : 56'h0; // @[DivSqrtRecFN_small.scala 342:12]
  assign _GEN_17 = {{1'd0}, _T_78}; // @[DivSqrtRecFN_small.scala 341:57]
  assign _T_87 = _GEN_17 | _T_86; // @[DivSqrtRecFN_small.scala 341:57]
  assign _T_89 = {rem_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 348:29]
  assign _T_90 = inReady ? 56'h0 : _T_89; // @[DivSqrtRecFN_small.scala 348:12]
  assign rem = _T_87 | _T_90; // @[DivSqrtRecFN_small.scala 347:11]
  assign bitMask = cycleNum[55:2]; // @[DivSqrtRecFN_small.scala 349:27]
  assign _T_92 = inReady & ~io_sqrtOp; // @[DivSqrtRecFN_small.scala 351:21]
  assign _T_93 = {io_b_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 351:47]
  assign _T_94 = _T_92 ? _T_93 : 55'h0; // @[DivSqrtRecFN_small.scala 351:12]
  assign _T_95 = inReady & evenSqrt_S; // @[DivSqrtRecFN_small.scala 352:21]
  assign _T_96 = _T_95 ? 54'h20000000000000 : 54'h0; // @[DivSqrtRecFN_small.scala 352:12]
  assign _GEN_18 = {{1'd0}, _T_96}; // @[DivSqrtRecFN_small.scala 351:73]
  assign _T_97 = _T_94 | _GEN_18; // @[DivSqrtRecFN_small.scala 351:73]
  assign _T_99 = _T_79 ? 55'h50000000000000 : 55'h0; // @[DivSqrtRecFN_small.scala 353:12]
  assign _T_100 = _T_97 | _T_99; // @[DivSqrtRecFN_small.scala 352:73]
  assign _T_103 = ~inReady & ~sqrtOp_Z; // @[DivSqrtRecFN_small.scala 354:23]
  assign _T_104 = {1'h1,fractB_Z}; // @[Cat.scala 29:58]
  assign _T_105 = {_T_104, 1'h0}; // @[DivSqrtRecFN_small.scala 354:56]
  assign _T_106 = _T_103 ? _T_105 : 54'h0; // @[DivSqrtRecFN_small.scala 354:12]
  assign _GEN_19 = {{1'd0}, _T_106}; // @[DivSqrtRecFN_small.scala 353:73]
  assign _T_107 = _T_100 | _GEN_19; // @[DivSqrtRecFN_small.scala 353:73]
  assign _T_109 = ~inReady & sqrtOp_Z; // @[DivSqrtRecFN_small.scala 355:23]
  assign _T_110 = {sigX_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 355:44]
  assign _GEN_20 = {{2'd0}, bitMask}; // @[DivSqrtRecFN_small.scala 355:48]
  assign _T_111 = _T_110 | _GEN_20; // @[DivSqrtRecFN_small.scala 355:48]
  assign _T_112 = _T_109 ? _T_111 : 56'h0; // @[DivSqrtRecFN_small.scala 355:12]
  assign _GEN_21 = {{1'd0}, _T_107}; // @[DivSqrtRecFN_small.scala 354:73]
  assign trialTerm = _GEN_21 | _T_112; // @[DivSqrtRecFN_small.scala 354:73]
  assign _T_113 = {1'b0,$signed(rem)}; // @[DivSqrtRecFN_small.scala 356:24]
  assign _T_114 = {1'b0,$signed(trialTerm)}; // @[DivSqrtRecFN_small.scala 356:41]
  assign trialRem = $signed(_T_113) - $signed(_T_114); // @[DivSqrtRecFN_small.scala 356:29]
  assign newBit = 57'sh0 <= $signed(trialRem); // @[DivSqrtRecFN_small.scala 357:23]
  assign _T_118 = idle | cycleNum[2]; // @[DivSqrtRecFN_small.scala 359:41]
  assign _T_120 = entering_normalCase | ~_T_118; // @[DivSqrtRecFN_small.scala 359:31]
  assign _T_121 = $signed(_T_113) - $signed(_T_114); // @[DivSqrtRecFN_small.scala 360:39]
  assign _T_122 = newBit ? _T_121 : {{1'd0}, rem}; // @[DivSqrtRecFN_small.scala 360:21]
  assign _GEN_10 = _T_120 ? _T_122 : {{2'd0}, rem_Z}; // @[DivSqrtRecFN_small.scala 359:58]
  assign _T_124 = ~inReady & newBit; // @[DivSqrtRecFN_small.scala 362:45]
  assign _T_125 = entering_normalCase | _T_124; // @[DivSqrtRecFN_small.scala 362:31]
  assign _T_126 = $signed(trialRem) != 57'sh0; // @[DivSqrtRecFN_small.scala 363:35]
  assign _T_129 = {newBit, 54'h0}; // @[DivSqrtRecFN_small.scala 365:47]
  assign _T_130 = _T_92 ? _T_129 : 55'h0; // @[DivSqrtRecFN_small.scala 365:16]
  assign _T_131 = inReady & io_sqrtOp; // @[DivSqrtRecFN_small.scala 366:25]
  assign _T_132 = _T_131 ? 54'h20000000000000 : 54'h0; // @[DivSqrtRecFN_small.scala 366:16]
  assign _GEN_22 = {{1'd0}, _T_132}; // @[DivSqrtRecFN_small.scala 365:71]
  assign _T_133 = _T_130 | _GEN_22; // @[DivSqrtRecFN_small.scala 365:71]
  assign _T_135 = {newBit, 52'h0}; // @[DivSqrtRecFN_small.scala 367:47]
  assign _T_136 = _T_79 ? _T_135 : 53'h0; // @[DivSqrtRecFN_small.scala 367:16]
  assign _GEN_23 = {{2'd0}, _T_136}; // @[DivSqrtRecFN_small.scala 366:71]
  assign _T_137 = _T_133 | _GEN_23; // @[DivSqrtRecFN_small.scala 366:71]
  assign _GEN_24 = {{1'd0}, bitMask}; // @[DivSqrtRecFN_small.scala 368:48]
  assign _T_139 = sigX_Z | _GEN_24; // @[DivSqrtRecFN_small.scala 368:48]
  assign _T_140 = inReady ? 55'h0 : _T_139; // @[DivSqrtRecFN_small.scala 368:16]
  assign _T_141 = _T_137 | _T_140; // @[DivSqrtRecFN_small.scala 367:71]
  assign _GEN_25 = {{55'd0}, notZeroRem_Z}; // @[DivSqrtRecFN_small.scala 385:35]
  assign io_inReady = idle | cycleNum[1]; // @[DivSqrtRecFN_small.scala 314:16]
  assign io_rawOutValid_div = cycleNum[1] & ~sqrtOp_Z; // @[DivSqrtRecFN_small.scala 375:25]
  assign io_rawOutValid_sqrt = cycleNum[1] & sqrtOp_Z; // @[DivSqrtRecFN_small.scala 376:25]
  assign io_roundingModeOut = roundingMode_Z; // @[DivSqrtRecFN_small.scala 377:25]
  assign io_invalidExc = majorExc_Z & isNaN_Z; // @[DivSqrtRecFN_small.scala 378:22]
  assign io_infiniteExc = majorExc_Z & ~isNaN_Z; // @[DivSqrtRecFN_small.scala 379:22]
  assign io_rawOut_isNaN = isNaN_Z; // @[DivSqrtRecFN_small.scala 380:22]
  assign io_rawOut_isInf = isInf_Z; // @[DivSqrtRecFN_small.scala 381:22]
  assign io_rawOut_isZero = isZero_Z; // @[DivSqrtRecFN_small.scala 382:22]
  assign io_rawOut_sign = sign_Z; // @[DivSqrtRecFN_small.scala 383:22]
  assign io_rawOut_sExp = sExp_Z; // @[DivSqrtRecFN_small.scala 384:22]
  assign io_rawOut_sig = _T_110 | _GEN_25; // @[DivSqrtRecFN_small.scala 385:22]
  assign DivSqrtRawFN_small_1_cov_read_addr = DivSqrtRawFN_small_1_state;
  assign DivSqrtRawFN_small_1_cov_read_data = DivSqrtRawFN_small_1_cov[DivSqrtRawFN_small_1_cov_read_addr]; // @[Coverage map for DivSqrtRawFN_small_1]
  assign DivSqrtRawFN_small_1_cov_write_data = 1'h1;
  assign DivSqrtRawFN_small_1_cov_write_addr = DivSqrtRawFN_small_1_state;
  assign DivSqrtRawFN_small_1_cov_write_mask = 1'h1;
  assign DivSqrtRawFN_small_1_cov_write_en = 1'h1;
  assign mux_cond_0 = _T_125;
  assign mux_cond_1 = newBit;
  assign mux_cond_2 = _T_63;
  assign mux_cond_3 = skipCycle2;
  assign sqrtOp_Z_shl = sqrtOp_Z;
  assign sqrtOp_Z_pad = {4'h0,sqrtOp_Z_shl};
  assign mux_cond_0_shl = {mux_cond_0, 1'h0};
  assign mux_cond_0_pad = {3'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 2'h0};
  assign mux_cond_1_pad = {2'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 3'h0};
  assign mux_cond_2_pad = {1'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 4'h0};
  assign mux_cond_3_pad = mux_cond_3_shl;
  assign DivSqrtRawFN_small_1_xor1 = sqrtOp_Z_pad ^ mux_cond_0_pad;
  assign DivSqrtRawFN_small_1_xor6 = mux_cond_2_pad ^ mux_cond_3_pad;
  assign DivSqrtRawFN_small_1_xor2 = mux_cond_1_pad ^ DivSqrtRawFN_small_1_xor6;
  assign DivSqrtRawFN_small_1_xor0 = DivSqrtRawFN_small_1_xor1 ^ DivSqrtRawFN_small_1_xor2;
  assign io_covSum = DivSqrtRawFN_small_1_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  cycleNum = _RAND_0[55:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  majorExc_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isNaN_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  isInf_Z = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  isZero_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sign_Z = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sExp_Z = _RAND_7[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  fractB_Z = _RAND_8[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  roundingMode_Z = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  rem_Z = _RAND_10[54:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  notZeroRem_Z = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sigX_Z = _RAND_12[54:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  DivSqrtRawFN_small_1_state = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    DivSqrtRawFN_small_1_cov[initvar] = _RAND_14[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  DivSqrtRawFN_small_1_covSum = _RAND_15[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      cycleNum <= 56'h0;
    end else if (reset) begin
      cycleNum <= 56'h1;
    end else if (_T_52) begin
      cycleNum <= _T_68;
    end
    if (metaReset) begin
      sqrtOp_Z <= 1'h0;
    end else if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (metaReset) begin
      majorExc_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        majorExc_Z <= _T_8;
      end else begin
        majorExc_Z <= _T_21;
      end
    end
    if (metaReset) begin
      isNaN_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isNaN_Z <= _T_22;
      end else begin
        isNaN_Z <= _T_24;
      end
    end
    if (metaReset) begin
      isInf_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isInf_Z <= io_a_isInf;
      end else begin
        isInf_Z <= _T_25;
      end
    end
    if (metaReset) begin
      isZero_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= io_a_isZero;
      end else begin
        isZero_Z <= _T_26;
      end
    end
    if (metaReset) begin
      sign_Z <= 1'h0;
    end else if (entering) begin
      sign_Z <= sign_S;
    end
    if (metaReset) begin
      sExp_Z <= 13'h0;
    end else if (entering_normalCase) begin
      if (io_sqrtOp) begin
        sExp_Z <= _T_70;
      end else begin
        sExp_Z <= sSatExpQuot_S_div;
      end
    end
    if (metaReset) begin
      fractB_Z <= 52'h0;
    end else if (_T_73) begin
      fractB_Z <= io_b_sig[51:0];
    end
    if (metaReset) begin
      roundingMode_Z <= 3'h0;
    end else if (entering_normalCase) begin
      roundingMode_Z <= io_roundingMode;
    end
    if (metaReset) begin
      rem_Z <= 55'h0;
    end else begin
      rem_Z <= _GEN_10[54:0];
    end
    if (metaReset) begin
      notZeroRem_Z <= 1'h0;
    end else if (_T_125) begin
      notZeroRem_Z <= _T_126;
    end
    if (metaReset) begin
      sigX_Z <= 55'h0;
    end else if (_T_125) begin
      sigX_Z <= _T_141;
    end
    DivSqrtRawFN_small_1_state <= DivSqrtRawFN_small_1_xor0;
    if (!(DivSqrtRawFN_small_1_cov_read_data)) begin
      DivSqrtRawFN_small_1_covSum <= DivSqrtRawFN_small_1_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(DivSqrtRawFN_small_1_cov_write_en & DivSqrtRawFN_small_1_cov_write_mask) begin
      DivSqrtRawFN_small_1_cov[DivSqrtRawFN_small_1_cov_write_addr] <= DivSqrtRawFN_small_1_cov_write_data; // @[Coverage map for DivSqrtRawFN_small_1]
    end
  end
endmodule
module RoundAnyRawFNToRecFN_6(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [55:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire  doShiftSigDown1; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire  _T_5; // @[primitives.scala 57:25]
  wire  _T_7; // @[primitives.scala 57:25]
  wire  _T_9; // @[primitives.scala 57:25]
  wire  _T_11; // @[primitives.scala 57:25]
  wire  _T_13; // @[primitives.scala 57:25]
  wire  _T_15; // @[primitives.scala 57:25]
  wire [5:0] _T_16; // @[primitives.scala 58:26]
  wire [64:0] _T_17; // @[primitives.scala 77:58]
  wire [31:0] _T_23; // @[Bitwise.scala 103:31]
  wire [31:0] _T_25; // @[Bitwise.scala 103:65]
  wire [31:0] _T_27; // @[Bitwise.scala 103:75]
  wire [31:0] _T_28; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_0; // @[Bitwise.scala 103:31]
  wire [31:0] _T_33; // @[Bitwise.scala 103:31]
  wire [31:0] _T_35; // @[Bitwise.scala 103:65]
  wire [31:0] _T_37; // @[Bitwise.scala 103:75]
  wire [31:0] _T_38; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [31:0] _T_43; // @[Bitwise.scala 103:31]
  wire [31:0] _T_45; // @[Bitwise.scala 103:65]
  wire [31:0] _T_47; // @[Bitwise.scala 103:75]
  wire [31:0] _T_48; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [31:0] _T_53; // @[Bitwise.scala 103:31]
  wire [31:0] _T_55; // @[Bitwise.scala 103:65]
  wire [31:0] _T_57; // @[Bitwise.scala 103:75]
  wire [31:0] _T_58; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_3; // @[Bitwise.scala 103:31]
  wire [31:0] _T_63; // @[Bitwise.scala 103:31]
  wire [31:0] _T_65; // @[Bitwise.scala 103:65]
  wire [31:0] _T_67; // @[Bitwise.scala 103:75]
  wire [31:0] _T_68; // @[Bitwise.scala 103:39]
  wire [15:0] _T_74; // @[Bitwise.scala 103:31]
  wire [15:0] _T_76; // @[Bitwise.scala 103:65]
  wire [15:0] _T_78; // @[Bitwise.scala 103:75]
  wire [15:0] _T_79; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_4; // @[Bitwise.scala 103:31]
  wire [15:0] _T_84; // @[Bitwise.scala 103:31]
  wire [15:0] _T_86; // @[Bitwise.scala 103:65]
  wire [15:0] _T_88; // @[Bitwise.scala 103:75]
  wire [15:0] _T_89; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_5; // @[Bitwise.scala 103:31]
  wire [15:0] _T_94; // @[Bitwise.scala 103:31]
  wire [15:0] _T_96; // @[Bitwise.scala 103:65]
  wire [15:0] _T_98; // @[Bitwise.scala 103:75]
  wire [15:0] _T_99; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_6; // @[Bitwise.scala 103:31]
  wire [15:0] _T_104; // @[Bitwise.scala 103:31]
  wire [15:0] _T_106; // @[Bitwise.scala 103:65]
  wire [15:0] _T_108; // @[Bitwise.scala 103:75]
  wire [15:0] _T_109; // @[Bitwise.scala 103:39]
  wire [50:0] _T_118; // @[Cat.scala 29:58]
  wire [50:0] _T_120; // @[primitives.scala 74:21]
  wire [50:0] _T_123; // @[primitives.scala 74:21]
  wire [50:0] _T_126; // @[primitives.scala 74:21]
  wire [50:0] _T_129; // @[primitives.scala 74:21]
  wire [53:0] _T_131; // @[Cat.scala 29:58]
  wire [2:0] _T_147; // @[Cat.scala 29:58]
  wire [2:0] _T_148; // @[primitives.scala 61:24]
  wire [2:0] _T_149; // @[primitives.scala 61:24]
  wire [2:0] _T_150; // @[primitives.scala 61:24]
  wire [2:0] _T_151; // @[primitives.scala 61:24]
  wire [53:0] _T_152; // @[primitives.scala 66:24]
  wire [53:0] _T_153; // @[primitives.scala 61:24]
  wire [53:0] _GEN_7; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [53:0] _T_154; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [55:0] _T_155; // @[Cat.scala 29:58]
  wire [55:0] _T_157; // @[Cat.scala 29:58]
  wire [55:0] _T_159; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [55:0] _T_160; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_161; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [55:0] _T_162; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_163; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  _T_164; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_165; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_166; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_167; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_168; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [55:0] _T_169; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [54:0] _T_171; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_172; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_174; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [54:0] _T_176; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [54:0] _T_178; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [55:0] _T_180; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_182; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [54:0] _T_184; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [54:0] _GEN_8; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _T_185; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _T_186; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_188; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [12:0] _GEN_9; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [13:0] _T_189; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [11:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [51:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _T_194; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  _T_199; // @[RoundAnyRawFNToRecFN.scala 201:16]
  wire  _T_201; // @[RoundAnyRawFNToRecFN.scala 203:30]
  wire  _T_203; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _T_204; // @[RoundAnyRawFNToRecFN.scala 203:49]
  wire  _T_206; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _T_207; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  _T_208; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire  _T_211; // @[RoundAnyRawFNToRecFN.scala 209:16]
  wire [1:0] _T_212; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _T_213; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _T_214; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _T_217; // @[RoundAnyRawFNToRecFN.scala 219:30]
  wire  _T_218; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _T_222; // @[RoundAnyRawFNToRecFN.scala 221:39]
  wire  _T_224; // @[RoundAnyRawFNToRecFN.scala 220:77]
  wire  _T_225; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _T_226; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _T_227; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _T_229; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 234:49]
  wire  _T_234; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _T_236; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _T_238; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _T_239; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _T_241; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _T_242; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [11:0] _T_243; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [11:0] _T_245; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [11:0] _T_247; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [11:0] _T_249; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [11:0] _T_250; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [11:0] _T_252; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [11:0] _T_253; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [11:0] _T_255; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [11:0] _T_256; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [11:0] _T_257; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [11:0] _T_258; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [11:0] _T_259; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [11:0] _T_260; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [11:0] _T_261; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [11:0] _T_262; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [11:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_263; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _T_264; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [51:0] _T_265; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [51:0] _T_266; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [51:0] _T_268; // @[Bitwise.scala 72:12]
  wire [51:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [12:0] _T_269; // @[Cat.scala 29:58]
  wire [1:0] _T_271; // @[Cat.scala 29:58]
  wire [2:0] _T_273; // @[Cat.scala 29:58]
  wire [29:0] RoundAnyRawFNToRecFN_6_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign doShiftSigDown1 = io_in_sig[55]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  assign _T_5 = ~io_in_sExp[11]; // @[primitives.scala 57:25]
  assign _T_7 = ~io_in_sExp[10]; // @[primitives.scala 57:25]
  assign _T_9 = ~io_in_sExp[9]; // @[primitives.scala 57:25]
  assign _T_11 = ~io_in_sExp[8]; // @[primitives.scala 57:25]
  assign _T_13 = ~io_in_sExp[7]; // @[primitives.scala 57:25]
  assign _T_15 = ~io_in_sExp[6]; // @[primitives.scala 57:25]
  assign _T_16 = ~io_in_sExp[5:0]; // @[primitives.scala 58:26]
  assign _T_17 = -65'sh10000000000000000 >>> _T_16; // @[primitives.scala 77:58]
  assign _T_23 = {{16'd0}, _T_17[44:29]}; // @[Bitwise.scala 103:31]
  assign _T_25 = {_T_17[28:13], 16'h0}; // @[Bitwise.scala 103:65]
  assign _T_27 = _T_25 & 32'hffff0000; // @[Bitwise.scala 103:75]
  assign _T_28 = _T_23 | _T_27; // @[Bitwise.scala 103:39]
  assign _GEN_0 = {{8'd0}, _T_28[31:8]}; // @[Bitwise.scala 103:31]
  assign _T_33 = _GEN_0 & 32'hff00ff; // @[Bitwise.scala 103:31]
  assign _T_35 = {_T_28[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_37 = _T_35 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  assign _T_38 = _T_33 | _T_37; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{4'd0}, _T_38[31:4]}; // @[Bitwise.scala 103:31]
  assign _T_43 = _GEN_1 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  assign _T_45 = {_T_38[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_47 = _T_45 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  assign _T_48 = _T_43 | _T_47; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{2'd0}, _T_48[31:2]}; // @[Bitwise.scala 103:31]
  assign _T_53 = _GEN_2 & 32'h33333333; // @[Bitwise.scala 103:31]
  assign _T_55 = {_T_48[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_57 = _T_55 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  assign _T_58 = _T_53 | _T_57; // @[Bitwise.scala 103:39]
  assign _GEN_3 = {{1'd0}, _T_58[31:1]}; // @[Bitwise.scala 103:31]
  assign _T_63 = _GEN_3 & 32'h55555555; // @[Bitwise.scala 103:31]
  assign _T_65 = {_T_58[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_67 = _T_65 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  assign _T_68 = _T_63 | _T_67; // @[Bitwise.scala 103:39]
  assign _T_74 = {{8'd0}, _T_17[60:53]}; // @[Bitwise.scala 103:31]
  assign _T_76 = {_T_17[52:45], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_78 = _T_76 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_79 = _T_74 | _T_78; // @[Bitwise.scala 103:39]
  assign _GEN_4 = {{4'd0}, _T_79[15:4]}; // @[Bitwise.scala 103:31]
  assign _T_84 = _GEN_4 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_86 = {_T_79[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_88 = _T_86 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_89 = _T_84 | _T_88; // @[Bitwise.scala 103:39]
  assign _GEN_5 = {{2'd0}, _T_89[15:2]}; // @[Bitwise.scala 103:31]
  assign _T_94 = _GEN_5 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_96 = {_T_89[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_98 = _T_96 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_99 = _T_94 | _T_98; // @[Bitwise.scala 103:39]
  assign _GEN_6 = {{1'd0}, _T_99[15:1]}; // @[Bitwise.scala 103:31]
  assign _T_104 = _GEN_6 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_106 = {_T_99[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_108 = _T_106 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_109 = _T_104 | _T_108; // @[Bitwise.scala 103:39]
  assign _T_118 = {_T_68,_T_109,_T_17[61],_T_17[62],_T_17[63]}; // @[Cat.scala 29:58]
  assign _T_120 = _T_15 ? 51'h0 : ~_T_118; // @[primitives.scala 74:21]
  assign _T_123 = _T_13 ? 51'h0 : _T_120[50:0]; // @[primitives.scala 74:21]
  assign _T_126 = _T_11 ? 51'h0 : _T_123[50:0]; // @[primitives.scala 74:21]
  assign _T_129 = _T_9 ? 51'h0 : _T_126[50:0]; // @[primitives.scala 74:21]
  assign _T_131 = {~_T_129,3'h7}; // @[Cat.scala 29:58]
  assign _T_147 = {_T_17[0],_T_17[1],_T_17[2]}; // @[Cat.scala 29:58]
  assign _T_148 = _T_15 ? _T_147 : 3'h0; // @[primitives.scala 61:24]
  assign _T_149 = _T_13 ? _T_148 : 3'h0; // @[primitives.scala 61:24]
  assign _T_150 = _T_11 ? _T_149 : 3'h0; // @[primitives.scala 61:24]
  assign _T_151 = _T_9 ? _T_150 : 3'h0; // @[primitives.scala 61:24]
  assign _T_152 = _T_7 ? _T_131 : {{51'd0}, _T_151}; // @[primitives.scala 66:24]
  assign _T_153 = _T_5 ? _T_152 : 54'h0; // @[primitives.scala 61:24]
  assign _GEN_7 = {{53'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_154 = _T_153 | _GEN_7; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_155 = {_T_154,2'h3}; // @[Cat.scala 29:58]
  assign _T_157 = {1'h0,_T_155[55:1]}; // @[Cat.scala 29:58]
  assign _T_159 = ~_T_157 & _T_155; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _T_160 = io_in_sig & _T_159; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_161 = |_T_160; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_162 = io_in_sig & _T_157; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_163 = |_T_162; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign _T_164 = _T_161 | _T_163; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_165 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_166 = _T_165 & _T_161; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_167 = roundMagUp & _T_164; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_168 = _T_166 | _T_167; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_169 = io_in_sig | _T_155; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_171 = _T_169[55:2] + 54'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_172 = roundingMode_near_even & _T_161; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_174 = _T_172 & ~_T_163; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_176 = _T_174 ? _T_155[55:1] : 55'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_178 = _T_171 & ~_T_176; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_180 = io_in_sig & ~_T_155; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_182 = roundingMode_odd & _T_164; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_184 = _T_182 ? _T_159[55:1] : 55'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_8 = {{1'd0}, _T_180[55:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_185 = _GEN_8 | _T_184; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_186 = _T_168 ? _T_178 : _T_185; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_188 = {1'b0,$signed(_T_186[54:53])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_9 = {{10{_T_188[2]}},_T_188}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_189 = $signed(io_in_sExp) + $signed(_GEN_9); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_189[11:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = doShiftSigDown1 ? _T_186[52:1] : _T_186[51:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  assign _T_194 = _T_189[13:10]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_T_194) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(_T_189) < 14'sh3ce; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign _T_199 = doShiftSigDown1 ? io_in_sig[2] : io_in_sig[1]; // @[RoundAnyRawFNToRecFN.scala 201:16]
  assign _T_201 = doShiftSigDown1 & io_in_sig[2]; // @[RoundAnyRawFNToRecFN.scala 203:30]
  assign _T_203 = |io_in_sig[1:0]; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign _T_204 = _T_201 | _T_203; // @[RoundAnyRawFNToRecFN.scala 203:49]
  assign _T_206 = _T_165 & _T_199; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _T_207 = roundMagUp & _T_204; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign _T_208 = _T_206 | _T_207; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign _T_211 = doShiftSigDown1 ? _T_186[54] : _T_186[53]; // @[RoundAnyRawFNToRecFN.scala 209:16]
  assign _T_212 = io_in_sExp[12:11]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _T_213 = $signed(_T_212) <= 2'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _T_214 = _T_164 & _T_213; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _T_217 = doShiftSigDown1 ? _T_155[3] : _T_155[2]; // @[RoundAnyRawFNToRecFN.scala 219:30]
  assign _T_218 = _T_214 & _T_217; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _T_222 = doShiftSigDown1 ? _T_155[4] : _T_155[3]; // @[RoundAnyRawFNToRecFN.scala 221:39]
  assign _T_224 = io_detectTininess & ~_T_222; // @[RoundAnyRawFNToRecFN.scala 220:77]
  assign _T_225 = _T_224 & _T_211; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _T_226 = _T_225 & _T_161; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _T_227 = _T_226 & _T_208; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _T_229 = _T_218 & ~_T_227; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _T_229; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | _T_164; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 234:49]
  assign _T_234 = ~isNaNOut & ~notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _T_234 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _T_236 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _T_236; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _T_165 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _T_238 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _T_239 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _T_238 & _T_239; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _T_241 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | _T_241; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _T_242 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _T_243 = _T_242 ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_245 = common_expOut & ~_T_243; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_247 = pegMinNonzeroMagOut ? 12'hc31 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _T_249 = _T_245 & ~_T_247; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _T_250 = pegMaxFiniteMagOut ? 12'h400 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _T_252 = _T_249 & ~_T_250; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _T_253 = notNaN_isInfOut ? 12'h200 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_255 = _T_252 & ~_T_253; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_256 = pegMinNonzeroMagOut ? 12'h3ce : 12'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _T_257 = _T_255 | _T_256; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _T_258 = pegMaxFiniteMagOut ? 12'hbff : 12'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _T_259 = _T_257 | _T_258; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _T_260 = notNaN_isInfOut ? 12'hc00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _T_261 = _T_259 | _T_260; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_262 = isNaNOut ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _T_261 | _T_262; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _T_263 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _T_264 = _T_263 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _T_265 = isNaNOut ? 52'h8000000000000 : 52'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _T_266 = _T_264 ? _T_265 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_268 = pegMaxFiniteMagOut ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  assign fractOut = _T_266 | _T_268; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign _T_269 = {signOut,expOut}; // @[Cat.scala 29:58]
  assign _T_271 = {underflow,inexact}; // @[Cat.scala 29:58]
  assign _T_273 = {io_invalidExc,io_infiniteExc,overflow}; // @[Cat.scala 29:58]
  assign io_out = {_T_269,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_273,_T_271}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_6_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_6_covSum;
  assign metaAssert = 1'h0;
endmodule
